module state_machine(	input logic Clk, Reset, Map, Battle);
endmodule