module register_file( input [15:0]

);

endmodule