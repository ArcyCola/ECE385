module datapath()

endmodule