module fakeramlmao (input clk, input[15:0] n, output pixelout );
always_ff @ (posedge clk)
begin
case (n)
0: pixelout<=1'b1;
1: pixelout<=1'b1;
2: pixelout<=1'b1;
3: pixelout<=1'b1;
4: pixelout<=1'b1;
5: pixelout<=1'b1;
6: pixelout<=1'b1;
7: pixelout<=1'b1;
8: pixelout<=1'b1;
9: pixelout<=1'b1;
10: pixelout<=1'b1;
11: pixelout<=1'b1;
12: pixelout<=1'b1;
13: pixelout<=1'b1;
14: pixelout<=1'b1;
15: pixelout<=1'b1;
16: pixelout<=1'b1;
17: pixelout<=1'b1;
18: pixelout<=1'b1;
19: pixelout<=1'b1;
20: pixelout<=1'b1;
21: pixelout<=1'b1;
22: pixelout<=1'b1;
23: pixelout<=1'b1;
24: pixelout<=1'b1;
25: pixelout<=1'b1;
26: pixelout<=1'b1;
27: pixelout<=1'b1;
28: pixelout<=1'b1;
29: pixelout<=1'b1;
30: pixelout<=1'b1;
31: pixelout<=1'b1;
32: pixelout<=1'b1;
33: pixelout<=1'b1;
34: pixelout<=1'b1;
35: pixelout<=1'b1;
36: pixelout<=1'b1;
37: pixelout<=1'b1;
38: pixelout<=1'b1;
39: pixelout<=1'b1;
40: pixelout<=1'b1;
41: pixelout<=1'b1;
42: pixelout<=1'b1;
43: pixelout<=1'b1;
44: pixelout<=1'b1;
45: pixelout<=1'b1;
46: pixelout<=1'b1;
47: pixelout<=1'b1;
48: pixelout<=1'b1;
49: pixelout<=1'b1;
50: pixelout<=1'b1;
51: pixelout<=1'b1;
52: pixelout<=1'b1;
53: pixelout<=1'b1;
54: pixelout<=1'b1;
55: pixelout<=1'b1;
56: pixelout<=1'b1;
57: pixelout<=1'b1;
58: pixelout<=1'b1;
59: pixelout<=1'b1;
60: pixelout<=1'b1;
61: pixelout<=1'b1;
62: pixelout<=1'b1;
63: pixelout<=1'b1;
64: pixelout<=1'b1;
65: pixelout<=1'b1;
66: pixelout<=1'b1;
67: pixelout<=1'b1;
68: pixelout<=1'b1;
69: pixelout<=1'b1;
70: pixelout<=1'b1;
71: pixelout<=1'b1;
72: pixelout<=1'b1;
73: pixelout<=1'b1;
74: pixelout<=1'b1;
75: pixelout<=1'b1;
76: pixelout<=1'b1;
77: pixelout<=1'b1;
78: pixelout<=1'b1;
79: pixelout<=1'b1;
80: pixelout<=1'b1;
81: pixelout<=1'b1;
82: pixelout<=1'b1;
83: pixelout<=1'b1;
84: pixelout<=1'b1;
85: pixelout<=1'b1;
86: pixelout<=1'b1;
87: pixelout<=1'b1;
88: pixelout<=1'b1;
89: pixelout<=1'b1;
90: pixelout<=1'b1;
91: pixelout<=1'b1;
92: pixelout<=1'b1;
93: pixelout<=1'b1;
94: pixelout<=1'b1;
95: pixelout<=1'b1;
96: pixelout<=1'b1;
97: pixelout<=1'b1;
98: pixelout<=1'b1;
99: pixelout<=1'b1;
100: pixelout<=1'b1;
101: pixelout<=1'b1;
102: pixelout<=1'b1;
103: pixelout<=1'b1;
104: pixelout<=1'b1;
105: pixelout<=1'b1;
106: pixelout<=1'b1;
107: pixelout<=1'b1;
108: pixelout<=1'b1;
109: pixelout<=1'b1;
110: pixelout<=1'b1;
111: pixelout<=1'b1;
112: pixelout<=1'b1;
113: pixelout<=1'b1;
114: pixelout<=1'b1;
115: pixelout<=1'b1;
116: pixelout<=1'b1;
117: pixelout<=1'b1;
118: pixelout<=1'b1;
119: pixelout<=1'b1;
120: pixelout<=1'b1;
121: pixelout<=1'b1;
122: pixelout<=1'b1;
123: pixelout<=1'b1;
124: pixelout<=1'b1;
125: pixelout<=1'b1;
126: pixelout<=1'b1;
127: pixelout<=1'b1;
128: pixelout<=1'b1;
129: pixelout<=1'b1;
130: pixelout<=1'b1;
131: pixelout<=1'b1;
132: pixelout<=1'b1;
133: pixelout<=1'b1;
134: pixelout<=1'b1;
135: pixelout<=1'b1;
136: pixelout<=1'b1;
137: pixelout<=1'b1;
138: pixelout<=1'b1;
139: pixelout<=1'b1;
140: pixelout<=1'b1;
141: pixelout<=1'b1;
142: pixelout<=1'b1;
143: pixelout<=1'b1;
144: pixelout<=1'b1;
145: pixelout<=1'b1;
146: pixelout<=1'b1;
147: pixelout<=1'b1;
148: pixelout<=1'b1;
149: pixelout<=1'b1;
150: pixelout<=1'b1;
151: pixelout<=1'b1;
152: pixelout<=1'b1;
153: pixelout<=1'b1;
154: pixelout<=1'b1;
155: pixelout<=1'b1;
156: pixelout<=1'b1;
157: pixelout<=1'b1;
158: pixelout<=1'b1;
159: pixelout<=1'b1;
160: pixelout<=1'b1;
161: pixelout<=1'b1;
162: pixelout<=1'b1;
163: pixelout<=1'b1;
164: pixelout<=1'b1;
165: pixelout<=1'b1;
166: pixelout<=1'b1;
167: pixelout<=1'b1;
168: pixelout<=1'b1;
169: pixelout<=1'b1;
170: pixelout<=1'b1;
171: pixelout<=1'b1;
172: pixelout<=1'b1;
173: pixelout<=1'b1;
174: pixelout<=1'b1;
175: pixelout<=1'b1;
176: pixelout<=1'b1;
177: pixelout<=1'b1;
178: pixelout<=1'b1;
179: pixelout<=1'b1;
180: pixelout<=1'b1;
181: pixelout<=1'b1;
182: pixelout<=1'b1;
183: pixelout<=1'b1;
184: pixelout<=1'b1;
185: pixelout<=1'b1;
186: pixelout<=1'b1;
187: pixelout<=1'b1;
188: pixelout<=1'b1;
189: pixelout<=1'b1;
190: pixelout<=1'b1;
191: pixelout<=1'b1;
192: pixelout<=1'b1;
193: pixelout<=1'b1;
194: pixelout<=1'b1;
195: pixelout<=1'b1;
196: pixelout<=1'b1;
197: pixelout<=1'b1;
198: pixelout<=1'b1;
199: pixelout<=1'b1;
200: pixelout<=1'b1;
201: pixelout<=1'b1;
202: pixelout<=1'b1;
203: pixelout<=1'b1;
204: pixelout<=1'b1;
205: pixelout<=1'b1;
206: pixelout<=1'b1;
207: pixelout<=1'b1;
208: pixelout<=1'b1;
209: pixelout<=1'b1;
210: pixelout<=1'b1;
211: pixelout<=1'b1;
212: pixelout<=1'b1;
213: pixelout<=1'b1;
214: pixelout<=1'b1;
215: pixelout<=1'b1;
216: pixelout<=1'b1;
217: pixelout<=1'b1;
218: pixelout<=1'b1;
219: pixelout<=1'b1;
220: pixelout<=1'b1;
221: pixelout<=1'b1;
222: pixelout<=1'b1;
223: pixelout<=1'b1;
224: pixelout<=1'b1;
225: pixelout<=1'b1;
226: pixelout<=1'b1;
227: pixelout<=1'b1;
228: pixelout<=1'b1;
229: pixelout<=1'b1;
230: pixelout<=1'b1;
231: pixelout<=1'b1;
232: pixelout<=1'b1;
233: pixelout<=1'b1;
234: pixelout<=1'b1;
235: pixelout<=1'b1;
236: pixelout<=1'b1;
237: pixelout<=1'b1;
238: pixelout<=1'b1;
239: pixelout<=1'b1;
240: pixelout<=1'b1;
241: pixelout<=1'b1;
242: pixelout<=1'b1;
243: pixelout<=1'b1;
244: pixelout<=1'b1;
245: pixelout<=1'b1;
246: pixelout<=1'b1;
247: pixelout<=1'b1;
248: pixelout<=1'b1;
249: pixelout<=1'b1;
250: pixelout<=1'b1;
251: pixelout<=1'b1;
252: pixelout<=1'b1;
253: pixelout<=1'b1;
254: pixelout<=1'b1;
255: pixelout<=1'b1;
256: pixelout<=1'b1;
257: pixelout<=1'b1;
258: pixelout<=1'b1;
259: pixelout<=1'b1;
260: pixelout<=1'b1;
261: pixelout<=1'b1;
262: pixelout<=1'b1;
263: pixelout<=1'b1;
264: pixelout<=1'b1;
265: pixelout<=1'b1;
266: pixelout<=1'b1;
267: pixelout<=1'b1;
268: pixelout<=1'b1;
269: pixelout<=1'b1;
270: pixelout<=1'b1;
271: pixelout<=1'b1;
272: pixelout<=1'b1;
273: pixelout<=1'b1;
274: pixelout<=1'b1;
275: pixelout<=1'b1;
276: pixelout<=1'b1;
277: pixelout<=1'b1;
278: pixelout<=1'b1;
279: pixelout<=1'b1;
280: pixelout<=1'b1;
281: pixelout<=1'b1;
282: pixelout<=1'b1;
283: pixelout<=1'b1;
284: pixelout<=1'b1;
285: pixelout<=1'b1;
286: pixelout<=1'b1;
287: pixelout<=1'b1;
288: pixelout<=1'b1;
289: pixelout<=1'b1;
290: pixelout<=1'b1;
291: pixelout<=1'b1;
292: pixelout<=1'b1;
293: pixelout<=1'b1;
294: pixelout<=1'b1;
295: pixelout<=1'b1;
296: pixelout<=1'b1;
297: pixelout<=1'b1;
298: pixelout<=1'b1;
299: pixelout<=1'b1;
300: pixelout<=1'b1;
301: pixelout<=1'b1;
302: pixelout<=1'b1;
303: pixelout<=1'b1;
304: pixelout<=1'b1;
305: pixelout<=1'b1;
306: pixelout<=1'b1;
307: pixelout<=1'b1;
308: pixelout<=1'b1;
309: pixelout<=1'b1;
310: pixelout<=1'b1;
311: pixelout<=1'b1;
312: pixelout<=1'b1;
313: pixelout<=1'b1;
314: pixelout<=1'b1;
315: pixelout<=1'b1;
316: pixelout<=1'b1;
317: pixelout<=1'b1;
318: pixelout<=1'b1;
319: pixelout<=1'b1;
320: pixelout<=1'b1;
321: pixelout<=1'b1;
322: pixelout<=1'b1;
323: pixelout<=1'b1;
324: pixelout<=1'b1;
325: pixelout<=1'b1;
326: pixelout<=1'b1;
327: pixelout<=1'b1;
328: pixelout<=1'b1;
329: pixelout<=1'b1;
330: pixelout<=1'b1;
331: pixelout<=1'b1;
332: pixelout<=1'b1;
333: pixelout<=1'b1;
334: pixelout<=1'b1;
335: pixelout<=1'b1;
336: pixelout<=1'b1;
337: pixelout<=1'b1;
338: pixelout<=1'b1;
339: pixelout<=1'b1;
340: pixelout<=1'b1;
341: pixelout<=1'b1;
342: pixelout<=1'b1;
343: pixelout<=1'b1;
344: pixelout<=1'b1;
345: pixelout<=1'b1;
346: pixelout<=1'b1;
347: pixelout<=1'b1;
348: pixelout<=1'b1;
349: pixelout<=1'b1;
350: pixelout<=1'b1;
351: pixelout<=1'b1;
352: pixelout<=1'b1;
353: pixelout<=1'b1;
354: pixelout<=1'b1;
355: pixelout<=1'b1;
356: pixelout<=1'b1;
357: pixelout<=1'b1;
358: pixelout<=1'b1;
359: pixelout<=1'b1;
360: pixelout<=1'b1;
361: pixelout<=1'b1;
362: pixelout<=1'b1;
363: pixelout<=1'b1;
364: pixelout<=1'b1;
365: pixelout<=1'b1;
366: pixelout<=1'b1;
367: pixelout<=1'b1;
368: pixelout<=1'b1;
369: pixelout<=1'b1;
370: pixelout<=1'b1;
371: pixelout<=1'b1;
372: pixelout<=1'b1;
373: pixelout<=1'b1;
374: pixelout<=1'b1;
375: pixelout<=1'b1;
376: pixelout<=1'b1;
377: pixelout<=1'b1;
378: pixelout<=1'b1;
379: pixelout<=1'b1;
380: pixelout<=1'b1;
381: pixelout<=1'b1;
382: pixelout<=1'b1;
383: pixelout<=1'b1;
384: pixelout<=1'b1;
385: pixelout<=1'b1;
386: pixelout<=1'b1;
387: pixelout<=1'b1;
388: pixelout<=1'b1;
389: pixelout<=1'b1;
390: pixelout<=1'b1;
391: pixelout<=1'b1;
392: pixelout<=1'b1;
393: pixelout<=1'b1;
394: pixelout<=1'b1;
395: pixelout<=1'b1;
396: pixelout<=1'b1;
397: pixelout<=1'b1;
398: pixelout<=1'b1;
399: pixelout<=1'b1;
400: pixelout<=1'b1;
401: pixelout<=1'b1;
402: pixelout<=1'b1;
403: pixelout<=1'b1;
404: pixelout<=1'b1;
405: pixelout<=1'b1;
406: pixelout<=1'b1;
407: pixelout<=1'b1;
408: pixelout<=1'b1;
409: pixelout<=1'b1;
410: pixelout<=1'b1;
411: pixelout<=1'b1;
412: pixelout<=1'b1;
413: pixelout<=1'b1;
414: pixelout<=1'b1;
415: pixelout<=1'b1;
416: pixelout<=1'b1;
417: pixelout<=1'b1;
418: pixelout<=1'b1;
419: pixelout<=1'b1;
420: pixelout<=1'b1;
421: pixelout<=1'b1;
422: pixelout<=1'b1;
423: pixelout<=1'b1;
424: pixelout<=1'b1;
425: pixelout<=1'b1;
426: pixelout<=1'b1;
427: pixelout<=1'b1;
428: pixelout<=1'b1;
429: pixelout<=1'b1;
430: pixelout<=1'b1;
431: pixelout<=1'b1;
432: pixelout<=1'b1;
433: pixelout<=1'b1;
434: pixelout<=1'b1;
435: pixelout<=1'b1;
436: pixelout<=1'b1;
437: pixelout<=1'b1;
438: pixelout<=1'b1;
439: pixelout<=1'b1;
440: pixelout<=1'b1;
441: pixelout<=1'b1;
442: pixelout<=1'b1;
443: pixelout<=1'b1;
444: pixelout<=1'b1;
445: pixelout<=1'b1;
446: pixelout<=1'b1;
447: pixelout<=1'b1;
448: pixelout<=1'b1;
449: pixelout<=1'b1;
450: pixelout<=1'b1;
451: pixelout<=1'b1;
452: pixelout<=1'b1;
453: pixelout<=1'b1;
454: pixelout<=1'b1;
455: pixelout<=1'b1;
456: pixelout<=1'b1;
457: pixelout<=1'b1;
458: pixelout<=1'b1;
459: pixelout<=1'b1;
460: pixelout<=1'b1;
461: pixelout<=1'b1;
462: pixelout<=1'b1;
463: pixelout<=1'b1;
464: pixelout<=1'b1;
465: pixelout<=1'b1;
466: pixelout<=1'b1;
467: pixelout<=1'b1;
468: pixelout<=1'b1;
469: pixelout<=1'b1;
470: pixelout<=1'b1;
471: pixelout<=1'b1;
472: pixelout<=1'b1;
473: pixelout<=1'b1;
474: pixelout<=1'b1;
475: pixelout<=1'b1;
476: pixelout<=1'b1;
477: pixelout<=1'b1;
478: pixelout<=1'b1;
479: pixelout<=1'b1;
480: pixelout<=1'b1;
481: pixelout<=1'b1;
482: pixelout<=1'b1;
483: pixelout<=1'b1;
484: pixelout<=1'b1;
485: pixelout<=1'b1;
486: pixelout<=1'b1;
487: pixelout<=1'b1;
488: pixelout<=1'b1;
489: pixelout<=1'b1;
490: pixelout<=1'b1;
491: pixelout<=1'b1;
492: pixelout<=1'b1;
493: pixelout<=1'b1;
494: pixelout<=1'b1;
495: pixelout<=1'b1;
496: pixelout<=1'b1;
497: pixelout<=1'b1;
498: pixelout<=1'b1;
499: pixelout<=1'b1;
500: pixelout<=1'b1;
501: pixelout<=1'b1;
502: pixelout<=1'b1;
503: pixelout<=1'b1;
504: pixelout<=1'b1;
505: pixelout<=1'b1;
506: pixelout<=1'b1;
507: pixelout<=1'b1;
508: pixelout<=1'b1;
509: pixelout<=1'b1;
510: pixelout<=1'b1;
511: pixelout<=1'b1;
512: pixelout<=1'b1;
513: pixelout<=1'b1;
514: pixelout<=1'b1;
515: pixelout<=1'b1;
516: pixelout<=1'b1;
517: pixelout<=1'b1;
518: pixelout<=1'b1;
519: pixelout<=1'b1;
520: pixelout<=1'b1;
521: pixelout<=1'b1;
522: pixelout<=1'b1;
523: pixelout<=1'b1;
524: pixelout<=1'b1;
525: pixelout<=1'b1;
526: pixelout<=1'b1;
527: pixelout<=1'b1;
528: pixelout<=1'b1;
529: pixelout<=1'b1;
530: pixelout<=1'b1;
531: pixelout<=1'b1;
532: pixelout<=1'b1;
533: pixelout<=1'b1;
534: pixelout<=1'b1;
535: pixelout<=1'b1;
536: pixelout<=1'b1;
537: pixelout<=1'b1;
538: pixelout<=1'b1;
539: pixelout<=1'b1;
540: pixelout<=1'b1;
541: pixelout<=1'b1;
542: pixelout<=1'b1;
543: pixelout<=1'b1;
544: pixelout<=1'b1;
545: pixelout<=1'b1;
546: pixelout<=1'b1;
547: pixelout<=1'b1;
548: pixelout<=1'b1;
549: pixelout<=1'b1;
550: pixelout<=1'b1;
551: pixelout<=1'b1;
552: pixelout<=1'b1;
553: pixelout<=1'b1;
554: pixelout<=1'b1;
555: pixelout<=1'b1;
556: pixelout<=1'b1;
557: pixelout<=1'b1;
558: pixelout<=1'b1;
559: pixelout<=1'b1;
560: pixelout<=1'b1;
561: pixelout<=1'b1;
562: pixelout<=1'b1;
563: pixelout<=1'b1;
564: pixelout<=1'b1;
565: pixelout<=1'b1;
566: pixelout<=1'b1;
567: pixelout<=1'b1;
568: pixelout<=1'b1;
569: pixelout<=1'b1;
570: pixelout<=1'b1;
571: pixelout<=1'b1;
572: pixelout<=1'b1;
573: pixelout<=1'b1;
574: pixelout<=1'b1;
575: pixelout<=1'b1;
576: pixelout<=1'b1;
577: pixelout<=1'b1;
578: pixelout<=1'b1;
579: pixelout<=1'b1;
580: pixelout<=1'b1;
581: pixelout<=1'b1;
582: pixelout<=1'b1;
583: pixelout<=1'b1;
584: pixelout<=1'b1;
585: pixelout<=1'b1;
586: pixelout<=1'b1;
587: pixelout<=1'b1;
588: pixelout<=1'b1;
589: pixelout<=1'b1;
590: pixelout<=1'b1;
591: pixelout<=1'b1;
592: pixelout<=1'b1;
593: pixelout<=1'b1;
594: pixelout<=1'b1;
595: pixelout<=1'b1;
596: pixelout<=1'b1;
597: pixelout<=1'b1;
598: pixelout<=1'b1;
599: pixelout<=1'b1;
600: pixelout<=1'b1;
601: pixelout<=1'b1;
602: pixelout<=1'b1;
603: pixelout<=1'b1;
604: pixelout<=1'b1;
605: pixelout<=1'b1;
606: pixelout<=1'b1;
607: pixelout<=1'b1;
608: pixelout<=1'b1;
609: pixelout<=1'b1;
610: pixelout<=1'b1;
611: pixelout<=1'b1;
612: pixelout<=1'b1;
613: pixelout<=1'b1;
614: pixelout<=1'b1;
615: pixelout<=1'b1;
616: pixelout<=1'b1;
617: pixelout<=1'b1;
618: pixelout<=1'b1;
619: pixelout<=1'b1;
620: pixelout<=1'b1;
621: pixelout<=1'b1;
622: pixelout<=1'b1;
623: pixelout<=1'b1;
624: pixelout<=1'b1;
625: pixelout<=1'b1;
626: pixelout<=1'b1;
627: pixelout<=1'b1;
628: pixelout<=1'b1;
629: pixelout<=1'b1;
630: pixelout<=1'b1;
631: pixelout<=1'b1;
632: pixelout<=1'b1;
633: pixelout<=1'b1;
634: pixelout<=1'b1;
635: pixelout<=1'b1;
636: pixelout<=1'b1;
637: pixelout<=1'b1;
638: pixelout<=1'b1;
639: pixelout<=1'b1;
640: pixelout<=1'b1;
641: pixelout<=1'b1;
642: pixelout<=1'b1;
643: pixelout<=1'b1;
644: pixelout<=1'b1;
645: pixelout<=1'b1;
646: pixelout<=1'b1;
647: pixelout<=1'b1;
648: pixelout<=1'b1;
649: pixelout<=1'b1;
650: pixelout<=1'b1;
651: pixelout<=1'b1;
652: pixelout<=1'b1;
653: pixelout<=1'b1;
654: pixelout<=1'b1;
655: pixelout<=1'b1;
656: pixelout<=1'b1;
657: pixelout<=1'b1;
658: pixelout<=1'b1;
659: pixelout<=1'b1;
660: pixelout<=1'b1;
661: pixelout<=1'b1;
662: pixelout<=1'b1;
663: pixelout<=1'b1;
664: pixelout<=1'b1;
665: pixelout<=1'b1;
666: pixelout<=1'b1;
667: pixelout<=1'b1;
668: pixelout<=1'b1;
669: pixelout<=1'b1;
670: pixelout<=1'b1;
671: pixelout<=1'b1;
672: pixelout<=1'b1;
673: pixelout<=1'b1;
674: pixelout<=1'b1;
675: pixelout<=1'b1;
676: pixelout<=1'b1;
677: pixelout<=1'b1;
678: pixelout<=1'b1;
679: pixelout<=1'b1;
680: pixelout<=1'b1;
681: pixelout<=1'b1;
682: pixelout<=1'b1;
683: pixelout<=1'b1;
684: pixelout<=1'b1;
685: pixelout<=1'b1;
686: pixelout<=1'b1;
687: pixelout<=1'b1;
688: pixelout<=1'b1;
689: pixelout<=1'b1;
690: pixelout<=1'b1;
691: pixelout<=1'b1;
692: pixelout<=1'b1;
693: pixelout<=1'b1;
694: pixelout<=1'b1;
695: pixelout<=1'b1;
696: pixelout<=1'b1;
697: pixelout<=1'b1;
698: pixelout<=1'b1;
699: pixelout<=1'b1;
700: pixelout<=1'b1;
701: pixelout<=1'b1;
702: pixelout<=1'b1;
703: pixelout<=1'b1;
704: pixelout<=1'b1;
705: pixelout<=1'b1;
706: pixelout<=1'b1;
707: pixelout<=1'b1;
708: pixelout<=1'b1;
709: pixelout<=1'b1;
710: pixelout<=1'b1;
711: pixelout<=1'b1;
712: pixelout<=1'b1;
713: pixelout<=1'b1;
714: pixelout<=1'b1;
715: pixelout<=1'b1;
716: pixelout<=1'b1;
717: pixelout<=1'b1;
718: pixelout<=1'b1;
719: pixelout<=1'b1;
720: pixelout<=1'b1;
721: pixelout<=1'b1;
722: pixelout<=1'b1;
723: pixelout<=1'b1;
724: pixelout<=1'b1;
725: pixelout<=1'b1;
726: pixelout<=1'b1;
727: pixelout<=1'b1;
728: pixelout<=1'b1;
729: pixelout<=1'b1;
730: pixelout<=1'b1;
731: pixelout<=1'b1;
732: pixelout<=1'b1;
733: pixelout<=1'b1;
734: pixelout<=1'b1;
735: pixelout<=1'b1;
736: pixelout<=1'b1;
737: pixelout<=1'b1;
738: pixelout<=1'b1;
739: pixelout<=1'b1;
740: pixelout<=1'b1;
741: pixelout<=1'b1;
742: pixelout<=1'b1;
743: pixelout<=1'b1;
744: pixelout<=1'b1;
745: pixelout<=1'b1;
746: pixelout<=1'b1;
747: pixelout<=1'b1;
748: pixelout<=1'b1;
749: pixelout<=1'b1;
750: pixelout<=1'b1;
751: pixelout<=1'b1;
752: pixelout<=1'b1;
753: pixelout<=1'b1;
754: pixelout<=1'b1;
755: pixelout<=1'b1;
756: pixelout<=1'b1;
757: pixelout<=1'b1;
758: pixelout<=1'b1;
759: pixelout<=1'b1;
760: pixelout<=1'b1;
761: pixelout<=1'b1;
762: pixelout<=1'b1;
763: pixelout<=1'b1;
764: pixelout<=1'b1;
765: pixelout<=1'b1;
766: pixelout<=1'b1;
767: pixelout<=1'b1;
768: pixelout<=1'b1;
769: pixelout<=1'b1;
770: pixelout<=1'b1;
771: pixelout<=1'b1;
772: pixelout<=1'b1;
773: pixelout<=1'b1;
774: pixelout<=1'b1;
775: pixelout<=1'b1;
776: pixelout<=1'b1;
777: pixelout<=1'b1;
778: pixelout<=1'b1;
779: pixelout<=1'b1;
780: pixelout<=1'b1;
781: pixelout<=1'b1;
782: pixelout<=1'b1;
783: pixelout<=1'b1;
784: pixelout<=1'b1;
785: pixelout<=1'b1;
786: pixelout<=1'b1;
787: pixelout<=1'b1;
788: pixelout<=1'b1;
789: pixelout<=1'b1;
790: pixelout<=1'b1;
791: pixelout<=1'b1;
792: pixelout<=1'b1;
793: pixelout<=1'b1;
794: pixelout<=1'b1;
795: pixelout<=1'b1;
796: pixelout<=1'b1;
797: pixelout<=1'b1;
798: pixelout<=1'b1;
799: pixelout<=1'b1;
800: pixelout<=1'b1;
801: pixelout<=1'b1;
802: pixelout<=1'b1;
803: pixelout<=1'b1;
804: pixelout<=1'b1;
805: pixelout<=1'b1;
806: pixelout<=1'b1;
807: pixelout<=1'b1;
808: pixelout<=1'b1;
809: pixelout<=1'b1;
810: pixelout<=1'b1;
811: pixelout<=1'b1;
812: pixelout<=1'b1;
813: pixelout<=1'b1;
814: pixelout<=1'b1;
815: pixelout<=1'b1;
816: pixelout<=1'b1;
817: pixelout<=1'b1;
818: pixelout<=1'b1;
819: pixelout<=1'b1;
820: pixelout<=1'b1;
821: pixelout<=1'b1;
822: pixelout<=1'b1;
823: pixelout<=1'b1;
824: pixelout<=1'b1;
825: pixelout<=1'b1;
826: pixelout<=1'b1;
827: pixelout<=1'b1;
828: pixelout<=1'b1;
829: pixelout<=1'b1;
830: pixelout<=1'b1;
831: pixelout<=1'b1;
832: pixelout<=1'b1;
833: pixelout<=1'b1;
834: pixelout<=1'b1;
835: pixelout<=1'b1;
836: pixelout<=1'b1;
837: pixelout<=1'b1;
838: pixelout<=1'b1;
839: pixelout<=1'b1;
840: pixelout<=1'b1;
841: pixelout<=1'b1;
842: pixelout<=1'b1;
843: pixelout<=1'b1;
844: pixelout<=1'b1;
845: pixelout<=1'b1;
846: pixelout<=1'b1;
847: pixelout<=1'b1;
848: pixelout<=1'b1;
849: pixelout<=1'b1;
850: pixelout<=1'b1;
851: pixelout<=1'b1;
852: pixelout<=1'b1;
853: pixelout<=1'b1;
854: pixelout<=1'b1;
855: pixelout<=1'b1;
856: pixelout<=1'b1;
857: pixelout<=1'b1;
858: pixelout<=1'b1;
859: pixelout<=1'b1;
860: pixelout<=1'b1;
861: pixelout<=1'b1;
862: pixelout<=1'b1;
863: pixelout<=1'b1;
864: pixelout<=1'b1;
865: pixelout<=1'b1;
866: pixelout<=1'b1;
867: pixelout<=1'b1;
868: pixelout<=1'b1;
869: pixelout<=1'b1;
870: pixelout<=1'b1;
871: pixelout<=1'b1;
872: pixelout<=1'b1;
873: pixelout<=1'b1;
874: pixelout<=1'b1;
875: pixelout<=1'b1;
876: pixelout<=1'b1;
877: pixelout<=1'b1;
878: pixelout<=1'b1;
879: pixelout<=1'b1;
880: pixelout<=1'b1;
881: pixelout<=1'b1;
882: pixelout<=1'b1;
883: pixelout<=1'b1;
884: pixelout<=1'b1;
885: pixelout<=1'b1;
886: pixelout<=1'b1;
887: pixelout<=1'b1;
888: pixelout<=1'b1;
889: pixelout<=1'b1;
890: pixelout<=1'b1;
891: pixelout<=1'b1;
892: pixelout<=1'b1;
893: pixelout<=1'b1;
894: pixelout<=1'b1;
895: pixelout<=1'b1;
896: pixelout<=1'b1;
897: pixelout<=1'b1;
898: pixelout<=1'b1;
899: pixelout<=1'b1;
900: pixelout<=1'b1;
901: pixelout<=1'b1;
902: pixelout<=1'b1;
903: pixelout<=1'b1;
904: pixelout<=1'b1;
905: pixelout<=1'b1;
906: pixelout<=1'b1;
907: pixelout<=1'b1;
908: pixelout<=1'b1;
909: pixelout<=1'b1;
910: pixelout<=1'b1;
911: pixelout<=1'b1;
912: pixelout<=1'b1;
913: pixelout<=1'b1;
914: pixelout<=1'b1;
915: pixelout<=1'b1;
916: pixelout<=1'b1;
917: pixelout<=1'b1;
918: pixelout<=1'b1;
919: pixelout<=1'b1;
920: pixelout<=1'b1;
921: pixelout<=1'b1;
922: pixelout<=1'b1;
923: pixelout<=1'b1;
924: pixelout<=1'b1;
925: pixelout<=1'b1;
926: pixelout<=1'b1;
927: pixelout<=1'b1;
928: pixelout<=1'b1;
929: pixelout<=1'b1;
930: pixelout<=1'b1;
931: pixelout<=1'b1;
932: pixelout<=1'b1;
933: pixelout<=1'b1;
934: pixelout<=1'b1;
935: pixelout<=1'b1;
936: pixelout<=1'b1;
937: pixelout<=1'b1;
938: pixelout<=1'b1;
939: pixelout<=1'b1;
940: pixelout<=1'b1;
941: pixelout<=1'b1;
942: pixelout<=1'b1;
943: pixelout<=1'b1;
944: pixelout<=1'b1;
945: pixelout<=1'b1;
946: pixelout<=1'b1;
947: pixelout<=1'b1;
948: pixelout<=1'b1;
949: pixelout<=1'b1;
950: pixelout<=1'b1;
951: pixelout<=1'b1;
952: pixelout<=1'b1;
953: pixelout<=1'b1;
954: pixelout<=1'b1;
955: pixelout<=1'b1;
956: pixelout<=1'b1;
957: pixelout<=1'b1;
958: pixelout<=1'b1;
959: pixelout<=1'b1;
960: pixelout<=1'b1;
961: pixelout<=1'b1;
962: pixelout<=1'b1;
963: pixelout<=1'b1;
964: pixelout<=1'b1;
965: pixelout<=1'b1;
966: pixelout<=1'b1;
967: pixelout<=1'b1;
968: pixelout<=1'b1;
969: pixelout<=1'b1;
970: pixelout<=1'b1;
971: pixelout<=1'b1;
972: pixelout<=1'b1;
973: pixelout<=1'b1;
974: pixelout<=1'b1;
975: pixelout<=1'b1;
976: pixelout<=1'b1;
977: pixelout<=1'b1;
978: pixelout<=1'b1;
979: pixelout<=1'b1;
980: pixelout<=1'b1;
981: pixelout<=1'b1;
982: pixelout<=1'b1;
983: pixelout<=1'b1;
984: pixelout<=1'b1;
985: pixelout<=1'b1;
986: pixelout<=1'b1;
987: pixelout<=1'b1;
988: pixelout<=1'b1;
989: pixelout<=1'b1;
990: pixelout<=1'b1;
991: pixelout<=1'b1;
992: pixelout<=1'b1;
993: pixelout<=1'b1;
994: pixelout<=1'b1;
995: pixelout<=1'b1;
996: pixelout<=1'b1;
997: pixelout<=1'b1;
998: pixelout<=1'b1;
999: pixelout<=1'b1;
1000: pixelout<=1'b1;
1001: pixelout<=1'b1;
1002: pixelout<=1'b1;
1003: pixelout<=1'b1;
1004: pixelout<=1'b1;
1005: pixelout<=1'b1;
1006: pixelout<=1'b1;
1007: pixelout<=1'b1;
1008: pixelout<=1'b1;
1009: pixelout<=1'b1;
1010: pixelout<=1'b1;
1011: pixelout<=1'b1;
1012: pixelout<=1'b1;
1013: pixelout<=1'b1;
1014: pixelout<=1'b1;
1015: pixelout<=1'b1;
1016: pixelout<=1'b1;
1017: pixelout<=1'b1;
1018: pixelout<=1'b1;
1019: pixelout<=1'b1;
1020: pixelout<=1'b1;
1021: pixelout<=1'b1;
1022: pixelout<=1'b1;
1023: pixelout<=1'b1;
1024: pixelout<=1'b1;
1025: pixelout<=1'b1;
1026: pixelout<=1'b1;
1027: pixelout<=1'b1;
1028: pixelout<=1'b1;
1029: pixelout<=1'b1;
1030: pixelout<=1'b1;
1031: pixelout<=1'b1;
1032: pixelout<=1'b1;
1033: pixelout<=1'b1;
1034: pixelout<=1'b1;
1035: pixelout<=1'b1;
1036: pixelout<=1'b1;
1037: pixelout<=1'b1;
1038: pixelout<=1'b1;
1039: pixelout<=1'b1;
1040: pixelout<=1'b1;
1041: pixelout<=1'b1;
1042: pixelout<=1'b1;
1043: pixelout<=1'b1;
1044: pixelout<=1'b1;
1045: pixelout<=1'b1;
1046: pixelout<=1'b1;
1047: pixelout<=1'b1;
1048: pixelout<=1'b1;
1049: pixelout<=1'b1;
1050: pixelout<=1'b1;
1051: pixelout<=1'b1;
1052: pixelout<=1'b1;
1053: pixelout<=1'b1;
1054: pixelout<=1'b1;
1055: pixelout<=1'b1;
1056: pixelout<=1'b1;
1057: pixelout<=1'b1;
1058: pixelout<=1'b1;
1059: pixelout<=1'b1;
1060: pixelout<=1'b1;
1061: pixelout<=1'b1;
1062: pixelout<=1'b1;
1063: pixelout<=1'b1;
1064: pixelout<=1'b1;
1065: pixelout<=1'b1;
1066: pixelout<=1'b1;
1067: pixelout<=1'b1;
1068: pixelout<=1'b1;
1069: pixelout<=1'b1;
1070: pixelout<=1'b1;
1071: pixelout<=1'b1;
1072: pixelout<=1'b1;
1073: pixelout<=1'b1;
1074: pixelout<=1'b1;
1075: pixelout<=1'b1;
1076: pixelout<=1'b1;
1077: pixelout<=1'b1;
1078: pixelout<=1'b1;
1079: pixelout<=1'b1;
1080: pixelout<=1'b1;
1081: pixelout<=1'b1;
1082: pixelout<=1'b1;
1083: pixelout<=1'b1;
1084: pixelout<=1'b1;
1085: pixelout<=1'b1;
1086: pixelout<=1'b1;
1087: pixelout<=1'b1;
1088: pixelout<=1'b1;
1089: pixelout<=1'b1;
1090: pixelout<=1'b1;
1091: pixelout<=1'b1;
1092: pixelout<=1'b1;
1093: pixelout<=1'b1;
1094: pixelout<=1'b1;
1095: pixelout<=1'b1;
1096: pixelout<=1'b1;
1097: pixelout<=1'b1;
1098: pixelout<=1'b1;
1099: pixelout<=1'b1;
1100: pixelout<=1'b1;
1101: pixelout<=1'b1;
1102: pixelout<=1'b1;
1103: pixelout<=1'b1;
1104: pixelout<=1'b1;
1105: pixelout<=1'b1;
1106: pixelout<=1'b1;
1107: pixelout<=1'b1;
1108: pixelout<=1'b1;
1109: pixelout<=1'b1;
1110: pixelout<=1'b1;
1111: pixelout<=1'b1;
1112: pixelout<=1'b1;
1113: pixelout<=1'b1;
1114: pixelout<=1'b1;
1115: pixelout<=1'b1;
1116: pixelout<=1'b1;
1117: pixelout<=1'b1;
1118: pixelout<=1'b1;
1119: pixelout<=1'b1;
1120: pixelout<=1'b1;
1121: pixelout<=1'b1;
1122: pixelout<=1'b1;
1123: pixelout<=1'b1;
1124: pixelout<=1'b1;
1125: pixelout<=1'b1;
1126: pixelout<=1'b1;
1127: pixelout<=1'b1;
1128: pixelout<=1'b1;
1129: pixelout<=1'b1;
1130: pixelout<=1'b1;
1131: pixelout<=1'b1;
1132: pixelout<=1'b1;
1133: pixelout<=1'b1;
1134: pixelout<=1'b1;
1135: pixelout<=1'b1;
1136: pixelout<=1'b1;
1137: pixelout<=1'b1;
1138: pixelout<=1'b1;
1139: pixelout<=1'b1;
1140: pixelout<=1'b1;
1141: pixelout<=1'b1;
1142: pixelout<=1'b1;
1143: pixelout<=1'b1;
1144: pixelout<=1'b1;
1145: pixelout<=1'b1;
1146: pixelout<=1'b1;
1147: pixelout<=1'b1;
1148: pixelout<=1'b1;
1149: pixelout<=1'b1;
1150: pixelout<=1'b1;
1151: pixelout<=1'b1;
1152: pixelout<=1'b1;
1153: pixelout<=1'b1;
1154: pixelout<=1'b1;
1155: pixelout<=1'b1;
1156: pixelout<=1'b1;
1157: pixelout<=1'b1;
1158: pixelout<=1'b1;
1159: pixelout<=1'b1;
1160: pixelout<=1'b1;
1161: pixelout<=1'b1;
1162: pixelout<=1'b1;
1163: pixelout<=1'b1;
1164: pixelout<=1'b1;
1165: pixelout<=1'b1;
1166: pixelout<=1'b1;
1167: pixelout<=1'b1;
1168: pixelout<=1'b1;
1169: pixelout<=1'b1;
1170: pixelout<=1'b1;
1171: pixelout<=1'b1;
1172: pixelout<=1'b1;
1173: pixelout<=1'b1;
1174: pixelout<=1'b1;
1175: pixelout<=1'b1;
1176: pixelout<=1'b1;
1177: pixelout<=1'b1;
1178: pixelout<=1'b1;
1179: pixelout<=1'b1;
1180: pixelout<=1'b1;
1181: pixelout<=1'b1;
1182: pixelout<=1'b1;
1183: pixelout<=1'b1;
1184: pixelout<=1'b1;
1185: pixelout<=1'b1;
1186: pixelout<=1'b1;
1187: pixelout<=1'b1;
1188: pixelout<=1'b1;
1189: pixelout<=1'b1;
1190: pixelout<=1'b1;
1191: pixelout<=1'b1;
1192: pixelout<=1'b1;
1193: pixelout<=1'b1;
1194: pixelout<=1'b1;
1195: pixelout<=1'b1;
1196: pixelout<=1'b1;
1197: pixelout<=1'b1;
1198: pixelout<=1'b1;
1199: pixelout<=1'b1;
1200: pixelout<=1'b1;
1201: pixelout<=1'b1;
1202: pixelout<=1'b1;
1203: pixelout<=1'b1;
1204: pixelout<=1'b1;
1205: pixelout<=1'b1;
1206: pixelout<=1'b1;
1207: pixelout<=1'b1;
1208: pixelout<=1'b1;
1209: pixelout<=1'b1;
1210: pixelout<=1'b1;
1211: pixelout<=1'b1;
1212: pixelout<=1'b1;
1213: pixelout<=1'b1;
1214: pixelout<=1'b1;
1215: pixelout<=1'b1;
1216: pixelout<=1'b1;
1217: pixelout<=1'b1;
1218: pixelout<=1'b1;
1219: pixelout<=1'b1;
1220: pixelout<=1'b1;
1221: pixelout<=1'b1;
1222: pixelout<=1'b1;
1223: pixelout<=1'b1;
1224: pixelout<=1'b1;
1225: pixelout<=1'b1;
1226: pixelout<=1'b1;
1227: pixelout<=1'b1;
1228: pixelout<=1'b1;
1229: pixelout<=1'b1;
1230: pixelout<=1'b1;
1231: pixelout<=1'b1;
1232: pixelout<=1'b1;
1233: pixelout<=1'b1;
1234: pixelout<=1'b1;
1235: pixelout<=1'b1;
1236: pixelout<=1'b1;
1237: pixelout<=1'b1;
1238: pixelout<=1'b1;
1239: pixelout<=1'b1;
1240: pixelout<=1'b1;
1241: pixelout<=1'b1;
1242: pixelout<=1'b1;
1243: pixelout<=1'b1;
1244: pixelout<=1'b1;
1245: pixelout<=1'b1;
1246: pixelout<=1'b1;
1247: pixelout<=1'b1;
1248: pixelout<=1'b1;
1249: pixelout<=1'b1;
1250: pixelout<=1'b1;
1251: pixelout<=1'b1;
1252: pixelout<=1'b1;
1253: pixelout<=1'b1;
1254: pixelout<=1'b1;
1255: pixelout<=1'b1;
1256: pixelout<=1'b1;
1257: pixelout<=1'b1;
1258: pixelout<=1'b1;
1259: pixelout<=1'b1;
1260: pixelout<=1'b1;
1261: pixelout<=1'b1;
1262: pixelout<=1'b1;
1263: pixelout<=1'b1;
1264: pixelout<=1'b1;
1265: pixelout<=1'b1;
1266: pixelout<=1'b1;
1267: pixelout<=1'b1;
1268: pixelout<=1'b1;
1269: pixelout<=1'b1;
1270: pixelout<=1'b1;
1271: pixelout<=1'b1;
1272: pixelout<=1'b1;
1273: pixelout<=1'b1;
1274: pixelout<=1'b1;
1275: pixelout<=1'b1;
1276: pixelout<=1'b1;
1277: pixelout<=1'b1;
1278: pixelout<=1'b1;
1279: pixelout<=1'b1;
1280: pixelout<=1'b1;
1281: pixelout<=1'b1;
1282: pixelout<=1'b1;
1283: pixelout<=1'b1;
1284: pixelout<=1'b1;
1285: pixelout<=1'b1;
1286: pixelout<=1'b1;
1287: pixelout<=1'b1;
1288: pixelout<=1'b1;
1289: pixelout<=1'b1;
1290: pixelout<=1'b1;
1291: pixelout<=1'b1;
1292: pixelout<=1'b1;
1293: pixelout<=1'b1;
1294: pixelout<=1'b1;
1295: pixelout<=1'b1;
1296: pixelout<=1'b1;
1297: pixelout<=1'b1;
1298: pixelout<=1'b1;
1299: pixelout<=1'b1;
1300: pixelout<=1'b1;
1301: pixelout<=1'b1;
1302: pixelout<=1'b1;
1303: pixelout<=1'b1;
1304: pixelout<=1'b1;
1305: pixelout<=1'b1;
1306: pixelout<=1'b1;
1307: pixelout<=1'b1;
1308: pixelout<=1'b1;
1309: pixelout<=1'b1;
1310: pixelout<=1'b1;
1311: pixelout<=1'b1;
1312: pixelout<=1'b1;
1313: pixelout<=1'b1;
1314: pixelout<=1'b1;
1315: pixelout<=1'b1;
1316: pixelout<=1'b1;
1317: pixelout<=1'b1;
1318: pixelout<=1'b1;
1319: pixelout<=1'b1;
1320: pixelout<=1'b1;
1321: pixelout<=1'b1;
1322: pixelout<=1'b1;
1323: pixelout<=1'b1;
1324: pixelout<=1'b1;
1325: pixelout<=1'b1;
1326: pixelout<=1'b1;
1327: pixelout<=1'b1;
1328: pixelout<=1'b1;
1329: pixelout<=1'b1;
1330: pixelout<=1'b1;
1331: pixelout<=1'b1;
1332: pixelout<=1'b1;
1333: pixelout<=1'b1;
1334: pixelout<=1'b1;
1335: pixelout<=1'b1;
1336: pixelout<=1'b1;
1337: pixelout<=1'b1;
1338: pixelout<=1'b1;
1339: pixelout<=1'b1;
1340: pixelout<=1'b1;
1341: pixelout<=1'b1;
1342: pixelout<=1'b1;
1343: pixelout<=1'b1;
1344: pixelout<=1'b1;
1345: pixelout<=1'b1;
1346: pixelout<=1'b1;
1347: pixelout<=1'b1;
1348: pixelout<=1'b1;
1349: pixelout<=1'b1;
1350: pixelout<=1'b1;
1351: pixelout<=1'b1;
1352: pixelout<=1'b1;
1353: pixelout<=1'b1;
1354: pixelout<=1'b1;
1355: pixelout<=1'b1;
1356: pixelout<=1'b1;
1357: pixelout<=1'b1;
1358: pixelout<=1'b1;
1359: pixelout<=1'b1;
1360: pixelout<=1'b1;
1361: pixelout<=1'b1;
1362: pixelout<=1'b1;
1363: pixelout<=1'b1;
1364: pixelout<=1'b1;
1365: pixelout<=1'b1;
1366: pixelout<=1'b1;
1367: pixelout<=1'b1;
1368: pixelout<=1'b1;
1369: pixelout<=1'b1;
1370: pixelout<=1'b1;
1371: pixelout<=1'b1;
1372: pixelout<=1'b1;
1373: pixelout<=1'b1;
1374: pixelout<=1'b1;
1375: pixelout<=1'b1;
1376: pixelout<=1'b1;
1377: pixelout<=1'b1;
1378: pixelout<=1'b1;
1379: pixelout<=1'b1;
1380: pixelout<=1'b1;
1381: pixelout<=1'b1;
1382: pixelout<=1'b1;
1383: pixelout<=1'b1;
1384: pixelout<=1'b1;
1385: pixelout<=1'b1;
1386: pixelout<=1'b1;
1387: pixelout<=1'b1;
1388: pixelout<=1'b1;
1389: pixelout<=1'b1;
1390: pixelout<=1'b1;
1391: pixelout<=1'b1;
1392: pixelout<=1'b1;
1393: pixelout<=1'b1;
1394: pixelout<=1'b1;
1395: pixelout<=1'b1;
1396: pixelout<=1'b1;
1397: pixelout<=1'b1;
1398: pixelout<=1'b1;
1399: pixelout<=1'b1;
1400: pixelout<=1'b1;
1401: pixelout<=1'b1;
1402: pixelout<=1'b1;
1403: pixelout<=1'b1;
1404: pixelout<=1'b1;
1405: pixelout<=1'b1;
1406: pixelout<=1'b1;
1407: pixelout<=1'b1;
1408: pixelout<=1'b1;
1409: pixelout<=1'b1;
1410: pixelout<=1'b1;
1411: pixelout<=1'b1;
1412: pixelout<=1'b1;
1413: pixelout<=1'b1;
1414: pixelout<=1'b1;
1415: pixelout<=1'b1;
1416: pixelout<=1'b1;
1417: pixelout<=1'b1;
1418: pixelout<=1'b1;
1419: pixelout<=1'b1;
1420: pixelout<=1'b1;
1421: pixelout<=1'b1;
1422: pixelout<=1'b1;
1423: pixelout<=1'b1;
1424: pixelout<=1'b1;
1425: pixelout<=1'b1;
1426: pixelout<=1'b1;
1427: pixelout<=1'b1;
1428: pixelout<=1'b1;
1429: pixelout<=1'b1;
1430: pixelout<=1'b1;
1431: pixelout<=1'b1;
1432: pixelout<=1'b1;
1433: pixelout<=1'b1;
1434: pixelout<=1'b1;
1435: pixelout<=1'b1;
1436: pixelout<=1'b1;
1437: pixelout<=1'b1;
1438: pixelout<=1'b1;
1439: pixelout<=1'b1;
1440: pixelout<=1'b1;
1441: pixelout<=1'b1;
1442: pixelout<=1'b1;
1443: pixelout<=1'b1;
1444: pixelout<=1'b1;
1445: pixelout<=1'b1;
1446: pixelout<=1'b1;
1447: pixelout<=1'b1;
1448: pixelout<=1'b1;
1449: pixelout<=1'b1;
1450: pixelout<=1'b1;
1451: pixelout<=1'b1;
1452: pixelout<=1'b1;
1453: pixelout<=1'b1;
1454: pixelout<=1'b1;
1455: pixelout<=1'b1;
1456: pixelout<=1'b1;
1457: pixelout<=1'b1;
1458: pixelout<=1'b1;
1459: pixelout<=1'b1;
1460: pixelout<=1'b1;
1461: pixelout<=1'b1;
1462: pixelout<=1'b1;
1463: pixelout<=1'b1;
1464: pixelout<=1'b1;
1465: pixelout<=1'b1;
1466: pixelout<=1'b1;
1467: pixelout<=1'b1;
1468: pixelout<=1'b1;
1469: pixelout<=1'b1;
1470: pixelout<=1'b1;
1471: pixelout<=1'b1;
1472: pixelout<=1'b1;
1473: pixelout<=1'b1;
1474: pixelout<=1'b1;
1475: pixelout<=1'b1;
1476: pixelout<=1'b1;
1477: pixelout<=1'b1;
1478: pixelout<=1'b1;
1479: pixelout<=1'b1;
1480: pixelout<=1'b1;
1481: pixelout<=1'b1;
1482: pixelout<=1'b1;
1483: pixelout<=1'b1;
1484: pixelout<=1'b1;
1485: pixelout<=1'b1;
1486: pixelout<=1'b1;
1487: pixelout<=1'b1;
1488: pixelout<=1'b1;
1489: pixelout<=1'b1;
1490: pixelout<=1'b1;
1491: pixelout<=1'b1;
1492: pixelout<=1'b1;
1493: pixelout<=1'b1;
1494: pixelout<=1'b1;
1495: pixelout<=1'b1;
1496: pixelout<=1'b1;
1497: pixelout<=1'b1;
1498: pixelout<=1'b1;
1499: pixelout<=1'b1;
1500: pixelout<=1'b1;
1501: pixelout<=1'b1;
1502: pixelout<=1'b1;
1503: pixelout<=1'b1;
1504: pixelout<=1'b1;
1505: pixelout<=1'b1;
1506: pixelout<=1'b1;
1507: pixelout<=1'b1;
1508: pixelout<=1'b1;
1509: pixelout<=1'b1;
1510: pixelout<=1'b1;
1511: pixelout<=1'b1;
1512: pixelout<=1'b1;
1513: pixelout<=1'b1;
1514: pixelout<=1'b1;
1515: pixelout<=1'b1;
1516: pixelout<=1'b1;
1517: pixelout<=1'b1;
1518: pixelout<=1'b1;
1519: pixelout<=1'b1;
1520: pixelout<=1'b1;
1521: pixelout<=1'b1;
1522: pixelout<=1'b1;
1523: pixelout<=1'b1;
1524: pixelout<=1'b1;
1525: pixelout<=1'b1;
1526: pixelout<=1'b1;
1527: pixelout<=1'b1;
1528: pixelout<=1'b1;
1529: pixelout<=1'b1;
1530: pixelout<=1'b1;
1531: pixelout<=1'b1;
1532: pixelout<=1'b1;
1533: pixelout<=1'b1;
1534: pixelout<=1'b1;
1535: pixelout<=1'b1;
1536: pixelout<=1'b1;
1537: pixelout<=1'b1;
1538: pixelout<=1'b1;
1539: pixelout<=1'b1;
1540: pixelout<=1'b1;
1541: pixelout<=1'b1;
1542: pixelout<=1'b1;
1543: pixelout<=1'b1;
1544: pixelout<=1'b1;
1545: pixelout<=1'b1;
1546: pixelout<=1'b1;
1547: pixelout<=1'b1;
1548: pixelout<=1'b1;
1549: pixelout<=1'b1;
1550: pixelout<=1'b1;
1551: pixelout<=1'b1;
1552: pixelout<=1'b1;
1553: pixelout<=1'b1;
1554: pixelout<=1'b1;
1555: pixelout<=1'b1;
1556: pixelout<=1'b1;
1557: pixelout<=1'b1;
1558: pixelout<=1'b1;
1559: pixelout<=1'b1;
1560: pixelout<=1'b1;
1561: pixelout<=1'b1;
1562: pixelout<=1'b1;
1563: pixelout<=1'b1;
1564: pixelout<=1'b1;
1565: pixelout<=1'b1;
1566: pixelout<=1'b1;
1567: pixelout<=1'b1;
1568: pixelout<=1'b1;
1569: pixelout<=1'b1;
1570: pixelout<=1'b1;
1571: pixelout<=1'b1;
1572: pixelout<=1'b1;
1573: pixelout<=1'b1;
1574: pixelout<=1'b1;
1575: pixelout<=1'b1;
1576: pixelout<=1'b1;
1577: pixelout<=1'b1;
1578: pixelout<=1'b1;
1579: pixelout<=1'b1;
1580: pixelout<=1'b1;
1581: pixelout<=1'b1;
1582: pixelout<=1'b1;
1583: pixelout<=1'b1;
1584: pixelout<=1'b1;
1585: pixelout<=1'b1;
1586: pixelout<=1'b1;
1587: pixelout<=1'b1;
1588: pixelout<=1'b1;
1589: pixelout<=1'b1;
1590: pixelout<=1'b1;
1591: pixelout<=1'b1;
1592: pixelout<=1'b1;
1593: pixelout<=1'b1;
1594: pixelout<=1'b1;
1595: pixelout<=1'b1;
1596: pixelout<=1'b1;
1597: pixelout<=1'b1;
1598: pixelout<=1'b1;
1599: pixelout<=1'b1;
1600: pixelout<=1'b1;
1601: pixelout<=1'b1;
1602: pixelout<=1'b1;
1603: pixelout<=1'b1;
1604: pixelout<=1'b1;
1605: pixelout<=1'b1;
1606: pixelout<=1'b1;
1607: pixelout<=1'b1;
1608: pixelout<=1'b1;
1609: pixelout<=1'b1;
1610: pixelout<=1'b1;
1611: pixelout<=1'b1;
1612: pixelout<=1'b1;
1613: pixelout<=1'b1;
1614: pixelout<=1'b1;
1615: pixelout<=1'b1;
1616: pixelout<=1'b1;
1617: pixelout<=1'b1;
1618: pixelout<=1'b1;
1619: pixelout<=1'b1;
1620: pixelout<=1'b1;
1621: pixelout<=1'b1;
1622: pixelout<=1'b1;
1623: pixelout<=1'b1;
1624: pixelout<=1'b1;
1625: pixelout<=1'b1;
1626: pixelout<=1'b1;
1627: pixelout<=1'b1;
1628: pixelout<=1'b1;
1629: pixelout<=1'b1;
1630: pixelout<=1'b1;
1631: pixelout<=1'b1;
1632: pixelout<=1'b1;
1633: pixelout<=1'b1;
1634: pixelout<=1'b1;
1635: pixelout<=1'b1;
1636: pixelout<=1'b1;
1637: pixelout<=1'b1;
1638: pixelout<=1'b1;
1639: pixelout<=1'b1;
1640: pixelout<=1'b1;
1641: pixelout<=1'b1;
1642: pixelout<=1'b1;
1643: pixelout<=1'b1;
1644: pixelout<=1'b1;
1645: pixelout<=1'b1;
1646: pixelout<=1'b1;
1647: pixelout<=1'b1;
1648: pixelout<=1'b1;
1649: pixelout<=1'b1;
1650: pixelout<=1'b1;
1651: pixelout<=1'b1;
1652: pixelout<=1'b1;
1653: pixelout<=1'b1;
1654: pixelout<=1'b1;
1655: pixelout<=1'b1;
1656: pixelout<=1'b1;
1657: pixelout<=1'b1;
1658: pixelout<=1'b1;
1659: pixelout<=1'b1;
1660: pixelout<=1'b1;
1661: pixelout<=1'b1;
1662: pixelout<=1'b1;
1663: pixelout<=1'b1;
1664: pixelout<=1'b1;
1665: pixelout<=1'b1;
1666: pixelout<=1'b1;
1667: pixelout<=1'b1;
1668: pixelout<=1'b1;
1669: pixelout<=1'b1;
1670: pixelout<=1'b1;
1671: pixelout<=1'b1;
1672: pixelout<=1'b1;
1673: pixelout<=1'b1;
1674: pixelout<=1'b1;
1675: pixelout<=1'b1;
1676: pixelout<=1'b1;
1677: pixelout<=1'b1;
1678: pixelout<=1'b1;
1679: pixelout<=1'b1;
1680: pixelout<=1'b1;
1681: pixelout<=1'b1;
1682: pixelout<=1'b1;
1683: pixelout<=1'b1;
1684: pixelout<=1'b1;
1685: pixelout<=1'b1;
1686: pixelout<=1'b1;
1687: pixelout<=1'b1;
1688: pixelout<=1'b1;
1689: pixelout<=1'b1;
1690: pixelout<=1'b1;
1691: pixelout<=1'b1;
1692: pixelout<=1'b1;
1693: pixelout<=1'b1;
1694: pixelout<=1'b1;
1695: pixelout<=1'b1;
1696: pixelout<=1'b1;
1697: pixelout<=1'b1;
1698: pixelout<=1'b1;
1699: pixelout<=1'b1;
1700: pixelout<=1'b1;
1701: pixelout<=1'b1;
1702: pixelout<=1'b1;
1703: pixelout<=1'b1;
1704: pixelout<=1'b1;
1705: pixelout<=1'b1;
1706: pixelout<=1'b1;
1707: pixelout<=1'b1;
1708: pixelout<=1'b1;
1709: pixelout<=1'b1;
1710: pixelout<=1'b1;
1711: pixelout<=1'b1;
1712: pixelout<=1'b1;
1713: pixelout<=1'b1;
1714: pixelout<=1'b1;
1715: pixelout<=1'b1;
1716: pixelout<=1'b1;
1717: pixelout<=1'b1;
1718: pixelout<=1'b1;
1719: pixelout<=1'b1;
1720: pixelout<=1'b1;
1721: pixelout<=1'b1;
1722: pixelout<=1'b1;
1723: pixelout<=1'b1;
1724: pixelout<=1'b1;
1725: pixelout<=1'b1;
1726: pixelout<=1'b1;
1727: pixelout<=1'b1;
1728: pixelout<=1'b1;
1729: pixelout<=1'b1;
1730: pixelout<=1'b1;
1731: pixelout<=1'b1;
1732: pixelout<=1'b1;
1733: pixelout<=1'b1;
1734: pixelout<=1'b1;
1735: pixelout<=1'b1;
1736: pixelout<=1'b1;
1737: pixelout<=1'b1;
1738: pixelout<=1'b1;
1739: pixelout<=1'b1;
1740: pixelout<=1'b1;
1741: pixelout<=1'b1;
1742: pixelout<=1'b1;
1743: pixelout<=1'b1;
1744: pixelout<=1'b1;
1745: pixelout<=1'b1;
1746: pixelout<=1'b1;
1747: pixelout<=1'b1;
1748: pixelout<=1'b1;
1749: pixelout<=1'b1;
1750: pixelout<=1'b1;
1751: pixelout<=1'b1;
1752: pixelout<=1'b1;
1753: pixelout<=1'b1;
1754: pixelout<=1'b1;
1755: pixelout<=1'b1;
1756: pixelout<=1'b1;
1757: pixelout<=1'b1;
1758: pixelout<=1'b1;
1759: pixelout<=1'b1;
1760: pixelout<=1'b1;
1761: pixelout<=1'b1;
1762: pixelout<=1'b1;
1763: pixelout<=1'b1;
1764: pixelout<=1'b1;
1765: pixelout<=1'b1;
1766: pixelout<=1'b1;
1767: pixelout<=1'b1;
1768: pixelout<=1'b1;
1769: pixelout<=1'b1;
1770: pixelout<=1'b1;
1771: pixelout<=1'b1;
1772: pixelout<=1'b1;
1773: pixelout<=1'b1;
1774: pixelout<=1'b1;
1775: pixelout<=1'b1;
1776: pixelout<=1'b1;
1777: pixelout<=1'b1;
1778: pixelout<=1'b1;
1779: pixelout<=1'b1;
1780: pixelout<=1'b1;
1781: pixelout<=1'b1;
1782: pixelout<=1'b1;
1783: pixelout<=1'b1;
1784: pixelout<=1'b1;
1785: pixelout<=1'b1;
1786: pixelout<=1'b1;
1787: pixelout<=1'b1;
1788: pixelout<=1'b1;
1789: pixelout<=1'b1;
1790: pixelout<=1'b1;
1791: pixelout<=1'b1;
1792: pixelout<=1'b1;
1793: pixelout<=1'b1;
1794: pixelout<=1'b1;
1795: pixelout<=1'b1;
1796: pixelout<=1'b1;
1797: pixelout<=1'b1;
1798: pixelout<=1'b1;
1799: pixelout<=1'b1;
1800: pixelout<=1'b1;
1801: pixelout<=1'b1;
1802: pixelout<=1'b1;
1803: pixelout<=1'b1;
1804: pixelout<=1'b1;
1805: pixelout<=1'b1;
1806: pixelout<=1'b1;
1807: pixelout<=1'b1;
1808: pixelout<=1'b1;
1809: pixelout<=1'b1;
1810: pixelout<=1'b1;
1811: pixelout<=1'b1;
1812: pixelout<=1'b1;
1813: pixelout<=1'b1;
1814: pixelout<=1'b1;
1815: pixelout<=1'b1;
1816: pixelout<=1'b1;
1817: pixelout<=1'b1;
1818: pixelout<=1'b1;
1819: pixelout<=1'b1;
1820: pixelout<=1'b1;
1821: pixelout<=1'b1;
1822: pixelout<=1'b1;
1823: pixelout<=1'b1;
1824: pixelout<=1'b1;
1825: pixelout<=1'b1;
1826: pixelout<=1'b1;
1827: pixelout<=1'b1;
1828: pixelout<=1'b1;
1829: pixelout<=1'b1;
1830: pixelout<=1'b1;
1831: pixelout<=1'b1;
1832: pixelout<=1'b1;
1833: pixelout<=1'b1;
1834: pixelout<=1'b1;
1835: pixelout<=1'b1;
1836: pixelout<=1'b1;
1837: pixelout<=1'b1;
1838: pixelout<=1'b1;
1839: pixelout<=1'b1;
1840: pixelout<=1'b1;
1841: pixelout<=1'b1;
1842: pixelout<=1'b1;
1843: pixelout<=1'b1;
1844: pixelout<=1'b1;
1845: pixelout<=1'b1;
1846: pixelout<=1'b1;
1847: pixelout<=1'b1;
1848: pixelout<=1'b1;
1849: pixelout<=1'b1;
1850: pixelout<=1'b1;
1851: pixelout<=1'b1;
1852: pixelout<=1'b1;
1853: pixelout<=1'b1;
1854: pixelout<=1'b1;
1855: pixelout<=1'b1;
1856: pixelout<=1'b1;
1857: pixelout<=1'b1;
1858: pixelout<=1'b1;
1859: pixelout<=1'b1;
1860: pixelout<=1'b1;
1861: pixelout<=1'b1;
1862: pixelout<=1'b1;
1863: pixelout<=1'b1;
1864: pixelout<=1'b1;
1865: pixelout<=1'b1;
1866: pixelout<=1'b1;
1867: pixelout<=1'b1;
1868: pixelout<=1'b1;
1869: pixelout<=1'b1;
1870: pixelout<=1'b1;
1871: pixelout<=1'b1;
1872: pixelout<=1'b1;
1873: pixelout<=1'b1;
1874: pixelout<=1'b1;
1875: pixelout<=1'b1;
1876: pixelout<=1'b1;
1877: pixelout<=1'b1;
1878: pixelout<=1'b1;
1879: pixelout<=1'b1;
1880: pixelout<=1'b1;
1881: pixelout<=1'b1;
1882: pixelout<=1'b1;
1883: pixelout<=1'b1;
1884: pixelout<=1'b1;
1885: pixelout<=1'b1;
1886: pixelout<=1'b1;
1887: pixelout<=1'b1;
1888: pixelout<=1'b1;
1889: pixelout<=1'b1;
1890: pixelout<=1'b1;
1891: pixelout<=1'b1;
1892: pixelout<=1'b1;
1893: pixelout<=1'b1;
1894: pixelout<=1'b1;
1895: pixelout<=1'b1;
1896: pixelout<=1'b1;
1897: pixelout<=1'b1;
1898: pixelout<=1'b1;
1899: pixelout<=1'b1;
1900: pixelout<=1'b1;
1901: pixelout<=1'b1;
1902: pixelout<=1'b1;
1903: pixelout<=1'b1;
1904: pixelout<=1'b1;
1905: pixelout<=1'b1;
1906: pixelout<=1'b1;
1907: pixelout<=1'b1;
1908: pixelout<=1'b1;
1909: pixelout<=1'b1;
1910: pixelout<=1'b1;
1911: pixelout<=1'b1;
1912: pixelout<=1'b1;
1913: pixelout<=1'b1;
1914: pixelout<=1'b1;
1915: pixelout<=1'b1;
1916: pixelout<=1'b1;
1917: pixelout<=1'b1;
1918: pixelout<=1'b1;
1919: pixelout<=1'b1;
1920: pixelout<=1'b1;
1921: pixelout<=1'b1;
1922: pixelout<=1'b1;
1923: pixelout<=1'b1;
1924: pixelout<=1'b1;
1925: pixelout<=1'b1;
1926: pixelout<=1'b1;
1927: pixelout<=1'b1;
1928: pixelout<=1'b1;
1929: pixelout<=1'b1;
1930: pixelout<=1'b1;
1931: pixelout<=1'b1;
1932: pixelout<=1'b1;
1933: pixelout<=1'b1;
1934: pixelout<=1'b1;
1935: pixelout<=1'b1;
1936: pixelout<=1'b1;
1937: pixelout<=1'b1;
1938: pixelout<=1'b1;
1939: pixelout<=1'b1;
1940: pixelout<=1'b1;
1941: pixelout<=1'b1;
1942: pixelout<=1'b1;
1943: pixelout<=1'b1;
1944: pixelout<=1'b1;
1945: pixelout<=1'b1;
1946: pixelout<=1'b1;
1947: pixelout<=1'b1;
1948: pixelout<=1'b1;
1949: pixelout<=1'b1;
1950: pixelout<=1'b1;
1951: pixelout<=1'b1;
1952: pixelout<=1'b1;
1953: pixelout<=1'b1;
1954: pixelout<=1'b1;
1955: pixelout<=1'b1;
1956: pixelout<=1'b1;
1957: pixelout<=1'b1;
1958: pixelout<=1'b1;
1959: pixelout<=1'b1;
1960: pixelout<=1'b1;
1961: pixelout<=1'b1;
1962: pixelout<=1'b1;
1963: pixelout<=1'b1;
1964: pixelout<=1'b1;
1965: pixelout<=1'b1;
1966: pixelout<=1'b1;
1967: pixelout<=1'b1;
1968: pixelout<=1'b1;
1969: pixelout<=1'b1;
1970: pixelout<=1'b1;
1971: pixelout<=1'b1;
1972: pixelout<=1'b1;
1973: pixelout<=1'b1;
1974: pixelout<=1'b1;
1975: pixelout<=1'b1;
1976: pixelout<=1'b1;
1977: pixelout<=1'b1;
1978: pixelout<=1'b1;
1979: pixelout<=1'b1;
1980: pixelout<=1'b1;
1981: pixelout<=1'b1;
1982: pixelout<=1'b1;
1983: pixelout<=1'b1;
1984: pixelout<=1'b1;
1985: pixelout<=1'b1;
1986: pixelout<=1'b1;
1987: pixelout<=1'b1;
1988: pixelout<=1'b1;
1989: pixelout<=1'b1;
1990: pixelout<=1'b1;
1991: pixelout<=1'b1;
1992: pixelout<=1'b1;
1993: pixelout<=1'b1;
1994: pixelout<=1'b1;
1995: pixelout<=1'b1;
1996: pixelout<=1'b1;
1997: pixelout<=1'b1;
1998: pixelout<=1'b1;
1999: pixelout<=1'b1;
2000: pixelout<=1'b1;
2001: pixelout<=1'b1;
2002: pixelout<=1'b1;
2003: pixelout<=1'b1;
2004: pixelout<=1'b1;
2005: pixelout<=1'b1;
2006: pixelout<=1'b1;
2007: pixelout<=1'b1;
2008: pixelout<=1'b1;
2009: pixelout<=1'b1;
2010: pixelout<=1'b1;
2011: pixelout<=1'b1;
2012: pixelout<=1'b1;
2013: pixelout<=1'b1;
2014: pixelout<=1'b1;
2015: pixelout<=1'b1;
2016: pixelout<=1'b1;
2017: pixelout<=1'b1;
2018: pixelout<=1'b1;
2019: pixelout<=1'b1;
2020: pixelout<=1'b1;
2021: pixelout<=1'b1;
2022: pixelout<=1'b1;
2023: pixelout<=1'b1;
2024: pixelout<=1'b1;
2025: pixelout<=1'b1;
2026: pixelout<=1'b1;
2027: pixelout<=1'b1;
2028: pixelout<=1'b1;
2029: pixelout<=1'b1;
2030: pixelout<=1'b1;
2031: pixelout<=1'b1;
2032: pixelout<=1'b1;
2033: pixelout<=1'b1;
2034: pixelout<=1'b1;
2035: pixelout<=1'b1;
2036: pixelout<=1'b1;
2037: pixelout<=1'b1;
2038: pixelout<=1'b1;
2039: pixelout<=1'b1;
2040: pixelout<=1'b1;
2041: pixelout<=1'b1;
2042: pixelout<=1'b1;
2043: pixelout<=1'b1;
2044: pixelout<=1'b1;
2045: pixelout<=1'b1;
2046: pixelout<=1'b1;
2047: pixelout<=1'b1;
2048: pixelout<=1'b1;
2049: pixelout<=1'b1;
2050: pixelout<=1'b1;
2051: pixelout<=1'b1;
2052: pixelout<=1'b1;
2053: pixelout<=1'b1;
2054: pixelout<=1'b1;
2055: pixelout<=1'b1;
2056: pixelout<=1'b1;
2057: pixelout<=1'b1;
2058: pixelout<=1'b1;
2059: pixelout<=1'b1;
2060: pixelout<=1'b1;
2061: pixelout<=1'b1;
2062: pixelout<=1'b1;
2063: pixelout<=1'b1;
2064: pixelout<=1'b1;
2065: pixelout<=1'b1;
2066: pixelout<=1'b1;
2067: pixelout<=1'b1;
2068: pixelout<=1'b1;
2069: pixelout<=1'b1;
2070: pixelout<=1'b1;
2071: pixelout<=1'b1;
2072: pixelout<=1'b1;
2073: pixelout<=1'b1;
2074: pixelout<=1'b1;
2075: pixelout<=1'b1;
2076: pixelout<=1'b1;
2077: pixelout<=1'b1;
2078: pixelout<=1'b1;
2079: pixelout<=1'b1;
2080: pixelout<=1'b1;
2081: pixelout<=1'b1;
2082: pixelout<=1'b1;
2083: pixelout<=1'b1;
2084: pixelout<=1'b1;
2085: pixelout<=1'b1;
2086: pixelout<=1'b1;
2087: pixelout<=1'b1;
2088: pixelout<=1'b1;
2089: pixelout<=1'b1;
2090: pixelout<=1'b1;
2091: pixelout<=1'b1;
2092: pixelout<=1'b1;
2093: pixelout<=1'b1;
2094: pixelout<=1'b1;
2095: pixelout<=1'b1;
2096: pixelout<=1'b1;
2097: pixelout<=1'b1;
2098: pixelout<=1'b1;
2099: pixelout<=1'b1;
2100: pixelout<=1'b1;
2101: pixelout<=1'b1;
2102: pixelout<=1'b1;
2103: pixelout<=1'b1;
2104: pixelout<=1'b1;
2105: pixelout<=1'b1;
2106: pixelout<=1'b1;
2107: pixelout<=1'b1;
2108: pixelout<=1'b1;
2109: pixelout<=1'b1;
2110: pixelout<=1'b1;
2111: pixelout<=1'b1;
2112: pixelout<=1'b1;
2113: pixelout<=1'b1;
2114: pixelout<=1'b1;
2115: pixelout<=1'b1;
2116: pixelout<=1'b1;
2117: pixelout<=1'b1;
2118: pixelout<=1'b1;
2119: pixelout<=1'b1;
2120: pixelout<=1'b1;
2121: pixelout<=1'b1;
2122: pixelout<=1'b1;
2123: pixelout<=1'b1;
2124: pixelout<=1'b1;
2125: pixelout<=1'b1;
2126: pixelout<=1'b1;
2127: pixelout<=1'b1;
2128: pixelout<=1'b1;
2129: pixelout<=1'b1;
2130: pixelout<=1'b1;
2131: pixelout<=1'b1;
2132: pixelout<=1'b1;
2133: pixelout<=1'b1;
2134: pixelout<=1'b1;
2135: pixelout<=1'b1;
2136: pixelout<=1'b1;
2137: pixelout<=1'b1;
2138: pixelout<=1'b1;
2139: pixelout<=1'b1;
2140: pixelout<=1'b1;
2141: pixelout<=1'b1;
2142: pixelout<=1'b1;
2143: pixelout<=1'b1;
2144: pixelout<=1'b1;
2145: pixelout<=1'b1;
2146: pixelout<=1'b1;
2147: pixelout<=1'b1;
2148: pixelout<=1'b1;
2149: pixelout<=1'b1;
2150: pixelout<=1'b1;
2151: pixelout<=1'b1;
2152: pixelout<=1'b1;
2153: pixelout<=1'b1;
2154: pixelout<=1'b1;
2155: pixelout<=1'b1;
2156: pixelout<=1'b1;
2157: pixelout<=1'b1;
2158: pixelout<=1'b1;
2159: pixelout<=1'b1;
2160: pixelout<=1'b1;
2161: pixelout<=1'b1;
2162: pixelout<=1'b1;
2163: pixelout<=1'b1;
2164: pixelout<=1'b1;
2165: pixelout<=1'b1;
2166: pixelout<=1'b1;
2167: pixelout<=1'b1;
2168: pixelout<=1'b1;
2169: pixelout<=1'b1;
2170: pixelout<=1'b1;
2171: pixelout<=1'b1;
2172: pixelout<=1'b1;
2173: pixelout<=1'b1;
2174: pixelout<=1'b1;
2175: pixelout<=1'b1;
2176: pixelout<=1'b1;
2177: pixelout<=1'b1;
2178: pixelout<=1'b1;
2179: pixelout<=1'b1;
2180: pixelout<=1'b1;
2181: pixelout<=1'b1;
2182: pixelout<=1'b1;
2183: pixelout<=1'b1;
2184: pixelout<=1'b1;
2185: pixelout<=1'b1;
2186: pixelout<=1'b1;
2187: pixelout<=1'b1;
2188: pixelout<=1'b1;
2189: pixelout<=1'b1;
2190: pixelout<=1'b1;
2191: pixelout<=1'b1;
2192: pixelout<=1'b1;
2193: pixelout<=1'b1;
2194: pixelout<=1'b1;
2195: pixelout<=1'b1;
2196: pixelout<=1'b1;
2197: pixelout<=1'b1;
2198: pixelout<=1'b1;
2199: pixelout<=1'b1;
2200: pixelout<=1'b1;
2201: pixelout<=1'b1;
2202: pixelout<=1'b1;
2203: pixelout<=1'b1;
2204: pixelout<=1'b1;
2205: pixelout<=1'b1;
2206: pixelout<=1'b1;
2207: pixelout<=1'b1;
2208: pixelout<=1'b1;
2209: pixelout<=1'b1;
2210: pixelout<=1'b1;
2211: pixelout<=1'b1;
2212: pixelout<=1'b1;
2213: pixelout<=1'b1;
2214: pixelout<=1'b1;
2215: pixelout<=1'b1;
2216: pixelout<=1'b1;
2217: pixelout<=1'b1;
2218: pixelout<=1'b1;
2219: pixelout<=1'b1;
2220: pixelout<=1'b1;
2221: pixelout<=1'b1;
2222: pixelout<=1'b1;
2223: pixelout<=1'b1;
2224: pixelout<=1'b1;
2225: pixelout<=1'b1;
2226: pixelout<=1'b1;
2227: pixelout<=1'b1;
2228: pixelout<=1'b1;
2229: pixelout<=1'b1;
2230: pixelout<=1'b1;
2231: pixelout<=1'b1;
2232: pixelout<=1'b1;
2233: pixelout<=1'b1;
2234: pixelout<=1'b1;
2235: pixelout<=1'b1;
2236: pixelout<=1'b1;
2237: pixelout<=1'b1;
2238: pixelout<=1'b1;
2239: pixelout<=1'b1;
2240: pixelout<=1'b1;
2241: pixelout<=1'b1;
2242: pixelout<=1'b1;
2243: pixelout<=1'b1;
2244: pixelout<=1'b1;
2245: pixelout<=1'b1;
2246: pixelout<=1'b1;
2247: pixelout<=1'b1;
2248: pixelout<=1'b1;
2249: pixelout<=1'b1;
2250: pixelout<=1'b1;
2251: pixelout<=1'b1;
2252: pixelout<=1'b1;
2253: pixelout<=1'b1;
2254: pixelout<=1'b1;
2255: pixelout<=1'b1;
2256: pixelout<=1'b1;
2257: pixelout<=1'b1;
2258: pixelout<=1'b1;
2259: pixelout<=1'b1;
2260: pixelout<=1'b1;
2261: pixelout<=1'b1;
2262: pixelout<=1'b1;
2263: pixelout<=1'b1;
2264: pixelout<=1'b1;
2265: pixelout<=1'b1;
2266: pixelout<=1'b1;
2267: pixelout<=1'b1;
2268: pixelout<=1'b1;
2269: pixelout<=1'b1;
2270: pixelout<=1'b1;
2271: pixelout<=1'b1;
2272: pixelout<=1'b1;
2273: pixelout<=1'b1;
2274: pixelout<=1'b1;
2275: pixelout<=1'b1;
2276: pixelout<=1'b1;
2277: pixelout<=1'b1;
2278: pixelout<=1'b1;
2279: pixelout<=1'b1;
2280: pixelout<=1'b1;
2281: pixelout<=1'b1;
2282: pixelout<=1'b1;
2283: pixelout<=1'b1;
2284: pixelout<=1'b1;
2285: pixelout<=1'b1;
2286: pixelout<=1'b1;
2287: pixelout<=1'b1;
2288: pixelout<=1'b1;
2289: pixelout<=1'b1;
2290: pixelout<=1'b1;
2291: pixelout<=1'b1;
2292: pixelout<=1'b1;
2293: pixelout<=1'b1;
2294: pixelout<=1'b1;
2295: pixelout<=1'b1;
2296: pixelout<=1'b1;
2297: pixelout<=1'b1;
2298: pixelout<=1'b1;
2299: pixelout<=1'b1;
2300: pixelout<=1'b1;
2301: pixelout<=1'b1;
2302: pixelout<=1'b1;
2303: pixelout<=1'b1;
2304: pixelout<=1'b1;
2305: pixelout<=1'b1;
2306: pixelout<=1'b1;
2307: pixelout<=1'b1;
2308: pixelout<=1'b1;
2309: pixelout<=1'b1;
2310: pixelout<=1'b1;
2311: pixelout<=1'b1;
2312: pixelout<=1'b1;
2313: pixelout<=1'b1;
2314: pixelout<=1'b1;
2315: pixelout<=1'b1;
2316: pixelout<=1'b1;
2317: pixelout<=1'b1;
2318: pixelout<=1'b1;
2319: pixelout<=1'b1;
2320: pixelout<=1'b1;
2321: pixelout<=1'b1;
2322: pixelout<=1'b1;
2323: pixelout<=1'b1;
2324: pixelout<=1'b1;
2325: pixelout<=1'b1;
2326: pixelout<=1'b1;
2327: pixelout<=1'b1;
2328: pixelout<=1'b1;
2329: pixelout<=1'b1;
2330: pixelout<=1'b1;
2331: pixelout<=1'b1;
2332: pixelout<=1'b1;
2333: pixelout<=1'b1;
2334: pixelout<=1'b1;
2335: pixelout<=1'b1;
2336: pixelout<=1'b1;
2337: pixelout<=1'b1;
2338: pixelout<=1'b1;
2339: pixelout<=1'b1;
2340: pixelout<=1'b1;
2341: pixelout<=1'b1;
2342: pixelout<=1'b1;
2343: pixelout<=1'b1;
2344: pixelout<=1'b1;
2345: pixelout<=1'b1;
2346: pixelout<=1'b1;
2347: pixelout<=1'b1;
2348: pixelout<=1'b1;
2349: pixelout<=1'b1;
2350: pixelout<=1'b1;
2351: pixelout<=1'b1;
2352: pixelout<=1'b1;
2353: pixelout<=1'b1;
2354: pixelout<=1'b1;
2355: pixelout<=1'b1;
2356: pixelout<=1'b1;
2357: pixelout<=1'b1;
2358: pixelout<=1'b1;
2359: pixelout<=1'b1;
2360: pixelout<=1'b1;
2361: pixelout<=1'b1;
2362: pixelout<=1'b1;
2363: pixelout<=1'b1;
2364: pixelout<=1'b1;
2365: pixelout<=1'b1;
2366: pixelout<=1'b1;
2367: pixelout<=1'b1;
2368: pixelout<=1'b1;
2369: pixelout<=1'b1;
2370: pixelout<=1'b1;
2371: pixelout<=1'b1;
2372: pixelout<=1'b1;
2373: pixelout<=1'b1;
2374: pixelout<=1'b1;
2375: pixelout<=1'b1;
2376: pixelout<=1'b1;
2377: pixelout<=1'b1;
2378: pixelout<=1'b1;
2379: pixelout<=1'b1;
2380: pixelout<=1'b1;
2381: pixelout<=1'b1;
2382: pixelout<=1'b1;
2383: pixelout<=1'b1;
2384: pixelout<=1'b1;
2385: pixelout<=1'b1;
2386: pixelout<=1'b1;
2387: pixelout<=1'b1;
2388: pixelout<=1'b1;
2389: pixelout<=1'b1;
2390: pixelout<=1'b1;
2391: pixelout<=1'b1;
2392: pixelout<=1'b1;
2393: pixelout<=1'b1;
2394: pixelout<=1'b1;
2395: pixelout<=1'b1;
2396: pixelout<=1'b1;
2397: pixelout<=1'b1;
2398: pixelout<=1'b1;
2399: pixelout<=1'b1;
2400: pixelout<=1'b1;
2401: pixelout<=1'b1;
2402: pixelout<=1'b1;
2403: pixelout<=1'b1;
2404: pixelout<=1'b1;
2405: pixelout<=1'b1;
2406: pixelout<=1'b1;
2407: pixelout<=1'b1;
2408: pixelout<=1'b1;
2409: pixelout<=1'b1;
2410: pixelout<=1'b1;
2411: pixelout<=1'b1;
2412: pixelout<=1'b1;
2413: pixelout<=1'b1;
2414: pixelout<=1'b1;
2415: pixelout<=1'b1;
2416: pixelout<=1'b1;
2417: pixelout<=1'b1;
2418: pixelout<=1'b1;
2419: pixelout<=1'b1;
2420: pixelout<=1'b1;
2421: pixelout<=1'b1;
2422: pixelout<=1'b1;
2423: pixelout<=1'b1;
2424: pixelout<=1'b1;
2425: pixelout<=1'b1;
2426: pixelout<=1'b1;
2427: pixelout<=1'b1;
2428: pixelout<=1'b1;
2429: pixelout<=1'b1;
2430: pixelout<=1'b1;
2431: pixelout<=1'b1;
2432: pixelout<=1'b1;
2433: pixelout<=1'b1;
2434: pixelout<=1'b1;
2435: pixelout<=1'b1;
2436: pixelout<=1'b1;
2437: pixelout<=1'b1;
2438: pixelout<=1'b1;
2439: pixelout<=1'b1;
2440: pixelout<=1'b1;
2441: pixelout<=1'b1;
2442: pixelout<=1'b1;
2443: pixelout<=1'b1;
2444: pixelout<=1'b1;
2445: pixelout<=1'b1;
2446: pixelout<=1'b1;
2447: pixelout<=1'b1;
2448: pixelout<=1'b1;
2449: pixelout<=1'b1;
2450: pixelout<=1'b0;
2451: pixelout<=1'b1;
2452: pixelout<=1'b1;
2453: pixelout<=1'b0;
2454: pixelout<=1'b1;
2455: pixelout<=1'b1;
2456: pixelout<=1'b1;
2457: pixelout<=1'b1;
2458: pixelout<=1'b1;
2459: pixelout<=1'b1;
2460: pixelout<=1'b1;
2461: pixelout<=1'b1;
2462: pixelout<=1'b1;
2463: pixelout<=1'b1;
2464: pixelout<=1'b1;
2465: pixelout<=1'b1;
2466: pixelout<=1'b1;
2467: pixelout<=1'b1;
2468: pixelout<=1'b1;
2469: pixelout<=1'b1;
2470: pixelout<=1'b1;
2471: pixelout<=1'b1;
2472: pixelout<=1'b1;
2473: pixelout<=1'b1;
2474: pixelout<=1'b1;
2475: pixelout<=1'b1;
2476: pixelout<=1'b1;
2477: pixelout<=1'b1;
2478: pixelout<=1'b1;
2479: pixelout<=1'b1;
2480: pixelout<=1'b1;
2481: pixelout<=1'b1;
2482: pixelout<=1'b1;
2483: pixelout<=1'b1;
2484: pixelout<=1'b1;
2485: pixelout<=1'b1;
2486: pixelout<=1'b1;
2487: pixelout<=1'b1;
2488: pixelout<=1'b1;
2489: pixelout<=1'b1;
2490: pixelout<=1'b1;
2491: pixelout<=1'b1;
2492: pixelout<=1'b1;
2493: pixelout<=1'b1;
2494: pixelout<=1'b1;
2495: pixelout<=1'b1;
2496: pixelout<=1'b1;
2497: pixelout<=1'b1;
2498: pixelout<=1'b1;
2499: pixelout<=1'b1;
2500: pixelout<=1'b1;
2501: pixelout<=1'b1;
2502: pixelout<=1'b1;
2503: pixelout<=1'b1;
2504: pixelout<=1'b1;
2505: pixelout<=1'b1;
2506: pixelout<=1'b1;
2507: pixelout<=1'b1;
2508: pixelout<=1'b1;
2509: pixelout<=1'b1;
2510: pixelout<=1'b1;
2511: pixelout<=1'b1;
2512: pixelout<=1'b1;
2513: pixelout<=1'b1;
2514: pixelout<=1'b1;
2515: pixelout<=1'b1;
2516: pixelout<=1'b1;
2517: pixelout<=1'b1;
2518: pixelout<=1'b1;
2519: pixelout<=1'b1;
2520: pixelout<=1'b1;
2521: pixelout<=1'b1;
2522: pixelout<=1'b1;
2523: pixelout<=1'b1;
2524: pixelout<=1'b1;
2525: pixelout<=1'b1;
2526: pixelout<=1'b1;
2527: pixelout<=1'b1;
2528: pixelout<=1'b1;
2529: pixelout<=1'b1;
2530: pixelout<=1'b1;
2531: pixelout<=1'b1;
2532: pixelout<=1'b1;
2533: pixelout<=1'b1;
2534: pixelout<=1'b1;
2535: pixelout<=1'b1;
2536: pixelout<=1'b1;
2537: pixelout<=1'b1;
2538: pixelout<=1'b1;
2539: pixelout<=1'b1;
2540: pixelout<=1'b1;
2541: pixelout<=1'b1;
2542: pixelout<=1'b1;
2543: pixelout<=1'b1;
2544: pixelout<=1'b1;
2545: pixelout<=1'b1;
2546: pixelout<=1'b1;
2547: pixelout<=1'b1;
2548: pixelout<=1'b1;
2549: pixelout<=1'b1;
2550: pixelout<=1'b1;
2551: pixelout<=1'b1;
2552: pixelout<=1'b1;
2553: pixelout<=1'b1;
2554: pixelout<=1'b1;
2555: pixelout<=1'b1;
2556: pixelout<=1'b1;
2557: pixelout<=1'b1;
2558: pixelout<=1'b1;
2559: pixelout<=1'b1;
2560: pixelout<=1'b1;
2561: pixelout<=1'b1;
2562: pixelout<=1'b1;
2563: pixelout<=1'b1;
2564: pixelout<=1'b1;
2565: pixelout<=1'b1;
2566: pixelout<=1'b1;
2567: pixelout<=1'b1;
2568: pixelout<=1'b1;
2569: pixelout<=1'b1;
2570: pixelout<=1'b1;
2571: pixelout<=1'b1;
2572: pixelout<=1'b1;
2573: pixelout<=1'b1;
2574: pixelout<=1'b1;
2575: pixelout<=1'b1;
2576: pixelout<=1'b1;
2577: pixelout<=1'b1;
2578: pixelout<=1'b1;
2579: pixelout<=1'b1;
2580: pixelout<=1'b1;
2581: pixelout<=1'b1;
2582: pixelout<=1'b1;
2583: pixelout<=1'b1;
2584: pixelout<=1'b1;
2585: pixelout<=1'b1;
2586: pixelout<=1'b1;
2587: pixelout<=1'b1;
2588: pixelout<=1'b1;
2589: pixelout<=1'b1;
2590: pixelout<=1'b1;
2591: pixelout<=1'b1;
2592: pixelout<=1'b1;
2593: pixelout<=1'b1;
2594: pixelout<=1'b1;
2595: pixelout<=1'b1;
2596: pixelout<=1'b1;
2597: pixelout<=1'b1;
2598: pixelout<=1'b1;
2599: pixelout<=1'b1;
2600: pixelout<=1'b1;
2601: pixelout<=1'b1;
2602: pixelout<=1'b1;
2603: pixelout<=1'b1;
2604: pixelout<=1'b1;
2605: pixelout<=1'b1;
2606: pixelout<=1'b1;
2607: pixelout<=1'b1;
2608: pixelout<=1'b1;
2609: pixelout<=1'b1;
2610: pixelout<=1'b1;
2611: pixelout<=1'b1;
2612: pixelout<=1'b1;
2613: pixelout<=1'b1;
2614: pixelout<=1'b1;
2615: pixelout<=1'b1;
2616: pixelout<=1'b1;
2617: pixelout<=1'b1;
2618: pixelout<=1'b1;
2619: pixelout<=1'b1;
2620: pixelout<=1'b1;
2621: pixelout<=1'b1;
2622: pixelout<=1'b1;
2623: pixelout<=1'b1;
2624: pixelout<=1'b1;
2625: pixelout<=1'b1;
2626: pixelout<=1'b1;
2627: pixelout<=1'b1;
2628: pixelout<=1'b1;
2629: pixelout<=1'b1;
2630: pixelout<=1'b1;
2631: pixelout<=1'b1;
2632: pixelout<=1'b1;
2633: pixelout<=1'b1;
2634: pixelout<=1'b1;
2635: pixelout<=1'b1;
2636: pixelout<=1'b1;
2637: pixelout<=1'b1;
2638: pixelout<=1'b1;
2639: pixelout<=1'b1;
2640: pixelout<=1'b1;
2641: pixelout<=1'b1;
2642: pixelout<=1'b1;
2643: pixelout<=1'b1;
2644: pixelout<=1'b1;
2645: pixelout<=1'b1;
2646: pixelout<=1'b1;
2647: pixelout<=1'b1;
2648: pixelout<=1'b1;
2649: pixelout<=1'b1;
2650: pixelout<=1'b1;
2651: pixelout<=1'b1;
2652: pixelout<=1'b1;
2653: pixelout<=1'b1;
2654: pixelout<=1'b1;
2655: pixelout<=1'b1;
2656: pixelout<=1'b1;
2657: pixelout<=1'b1;
2658: pixelout<=1'b1;
2659: pixelout<=1'b1;
2660: pixelout<=1'b1;
2661: pixelout<=1'b1;
2662: pixelout<=1'b1;
2663: pixelout<=1'b1;
2664: pixelout<=1'b1;
2665: pixelout<=1'b1;
2666: pixelout<=1'b1;
2667: pixelout<=1'b1;
2668: pixelout<=1'b1;
2669: pixelout<=1'b1;
2670: pixelout<=1'b1;
2671: pixelout<=1'b1;
2672: pixelout<=1'b1;
2673: pixelout<=1'b1;
2674: pixelout<=1'b1;
2675: pixelout<=1'b1;
2676: pixelout<=1'b1;
2677: pixelout<=1'b1;
2678: pixelout<=1'b1;
2679: pixelout<=1'b1;
2680: pixelout<=1'b1;
2681: pixelout<=1'b1;
2682: pixelout<=1'b1;
2683: pixelout<=1'b1;
2684: pixelout<=1'b1;
2685: pixelout<=1'b1;
2686: pixelout<=1'b1;
2687: pixelout<=1'b1;
2688: pixelout<=1'b1;
2689: pixelout<=1'b1;
2690: pixelout<=1'b0;
2691: pixelout<=1'b0;
2692: pixelout<=1'b1;
2693: pixelout<=1'b0;
2694: pixelout<=1'b0;
2695: pixelout<=1'b1;
2696: pixelout<=1'b1;
2697: pixelout<=1'b1;
2698: pixelout<=1'b1;
2699: pixelout<=1'b1;
2700: pixelout<=1'b1;
2701: pixelout<=1'b1;
2702: pixelout<=1'b1;
2703: pixelout<=1'b1;
2704: pixelout<=1'b1;
2705: pixelout<=1'b1;
2706: pixelout<=1'b1;
2707: pixelout<=1'b1;
2708: pixelout<=1'b1;
2709: pixelout<=1'b1;
2710: pixelout<=1'b1;
2711: pixelout<=1'b1;
2712: pixelout<=1'b1;
2713: pixelout<=1'b1;
2714: pixelout<=1'b1;
2715: pixelout<=1'b1;
2716: pixelout<=1'b1;
2717: pixelout<=1'b1;
2718: pixelout<=1'b1;
2719: pixelout<=1'b1;
2720: pixelout<=1'b1;
2721: pixelout<=1'b1;
2722: pixelout<=1'b1;
2723: pixelout<=1'b1;
2724: pixelout<=1'b1;
2725: pixelout<=1'b1;
2726: pixelout<=1'b1;
2727: pixelout<=1'b1;
2728: pixelout<=1'b1;
2729: pixelout<=1'b1;
2730: pixelout<=1'b1;
2731: pixelout<=1'b1;
2732: pixelout<=1'b1;
2733: pixelout<=1'b1;
2734: pixelout<=1'b1;
2735: pixelout<=1'b1;
2736: pixelout<=1'b1;
2737: pixelout<=1'b1;
2738: pixelout<=1'b1;
2739: pixelout<=1'b1;
2740: pixelout<=1'b1;
2741: pixelout<=1'b1;
2742: pixelout<=1'b0;
2743: pixelout<=1'b1;
2744: pixelout<=1'b1;
2745: pixelout<=1'b1;
2746: pixelout<=1'b1;
2747: pixelout<=1'b1;
2748: pixelout<=1'b1;
2749: pixelout<=1'b1;
2750: pixelout<=1'b1;
2751: pixelout<=1'b1;
2752: pixelout<=1'b1;
2753: pixelout<=1'b1;
2754: pixelout<=1'b1;
2755: pixelout<=1'b1;
2756: pixelout<=1'b1;
2757: pixelout<=1'b1;
2758: pixelout<=1'b1;
2759: pixelout<=1'b1;
2760: pixelout<=1'b1;
2761: pixelout<=1'b1;
2762: pixelout<=1'b1;
2763: pixelout<=1'b1;
2764: pixelout<=1'b1;
2765: pixelout<=1'b1;
2766: pixelout<=1'b1;
2767: pixelout<=1'b1;
2768: pixelout<=1'b1;
2769: pixelout<=1'b1;
2770: pixelout<=1'b1;
2771: pixelout<=1'b1;
2772: pixelout<=1'b1;
2773: pixelout<=1'b1;
2774: pixelout<=1'b1;
2775: pixelout<=1'b1;
2776: pixelout<=1'b1;
2777: pixelout<=1'b1;
2778: pixelout<=1'b1;
2779: pixelout<=1'b1;
2780: pixelout<=1'b1;
2781: pixelout<=1'b1;
2782: pixelout<=1'b1;
2783: pixelout<=1'b1;
2784: pixelout<=1'b1;
2785: pixelout<=1'b1;
2786: pixelout<=1'b1;
2787: pixelout<=1'b1;
2788: pixelout<=1'b1;
2789: pixelout<=1'b1;
2790: pixelout<=1'b1;
2791: pixelout<=1'b1;
2792: pixelout<=1'b1;
2793: pixelout<=1'b1;
2794: pixelout<=1'b1;
2795: pixelout<=1'b1;
2796: pixelout<=1'b1;
2797: pixelout<=1'b1;
2798: pixelout<=1'b1;
2799: pixelout<=1'b1;
2800: pixelout<=1'b1;
2801: pixelout<=1'b1;
2802: pixelout<=1'b1;
2803: pixelout<=1'b1;
2804: pixelout<=1'b1;
2805: pixelout<=1'b1;
2806: pixelout<=1'b1;
2807: pixelout<=1'b1;
2808: pixelout<=1'b1;
2809: pixelout<=1'b1;
2810: pixelout<=1'b1;
2811: pixelout<=1'b1;
2812: pixelout<=1'b1;
2813: pixelout<=1'b1;
2814: pixelout<=1'b1;
2815: pixelout<=1'b1;
2816: pixelout<=1'b1;
2817: pixelout<=1'b1;
2818: pixelout<=1'b1;
2819: pixelout<=1'b1;
2820: pixelout<=1'b1;
2821: pixelout<=1'b1;
2822: pixelout<=1'b1;
2823: pixelout<=1'b1;
2824: pixelout<=1'b1;
2825: pixelout<=1'b1;
2826: pixelout<=1'b1;
2827: pixelout<=1'b1;
2828: pixelout<=1'b1;
2829: pixelout<=1'b1;
2830: pixelout<=1'b1;
2831: pixelout<=1'b1;
2832: pixelout<=1'b1;
2833: pixelout<=1'b1;
2834: pixelout<=1'b1;
2835: pixelout<=1'b1;
2836: pixelout<=1'b1;
2837: pixelout<=1'b1;
2838: pixelout<=1'b1;
2839: pixelout<=1'b1;
2840: pixelout<=1'b1;
2841: pixelout<=1'b1;
2842: pixelout<=1'b1;
2843: pixelout<=1'b1;
2844: pixelout<=1'b1;
2845: pixelout<=1'b1;
2846: pixelout<=1'b1;
2847: pixelout<=1'b1;
2848: pixelout<=1'b1;
2849: pixelout<=1'b1;
2850: pixelout<=1'b1;
2851: pixelout<=1'b1;
2852: pixelout<=1'b1;
2853: pixelout<=1'b1;
2854: pixelout<=1'b1;
2855: pixelout<=1'b1;
2856: pixelout<=1'b1;
2857: pixelout<=1'b1;
2858: pixelout<=1'b1;
2859: pixelout<=1'b1;
2860: pixelout<=1'b1;
2861: pixelout<=1'b1;
2862: pixelout<=1'b1;
2863: pixelout<=1'b1;
2864: pixelout<=1'b1;
2865: pixelout<=1'b1;
2866: pixelout<=1'b1;
2867: pixelout<=1'b1;
2868: pixelout<=1'b1;
2869: pixelout<=1'b1;
2870: pixelout<=1'b1;
2871: pixelout<=1'b1;
2872: pixelout<=1'b1;
2873: pixelout<=1'b1;
2874: pixelout<=1'b1;
2875: pixelout<=1'b1;
2876: pixelout<=1'b1;
2877: pixelout<=1'b1;
2878: pixelout<=1'b1;
2879: pixelout<=1'b1;
2880: pixelout<=1'b1;
2881: pixelout<=1'b1;
2882: pixelout<=1'b1;
2883: pixelout<=1'b1;
2884: pixelout<=1'b1;
2885: pixelout<=1'b1;
2886: pixelout<=1'b1;
2887: pixelout<=1'b1;
2888: pixelout<=1'b1;
2889: pixelout<=1'b1;
2890: pixelout<=1'b1;
2891: pixelout<=1'b1;
2892: pixelout<=1'b1;
2893: pixelout<=1'b1;
2894: pixelout<=1'b1;
2895: pixelout<=1'b1;
2896: pixelout<=1'b1;
2897: pixelout<=1'b1;
2898: pixelout<=1'b1;
2899: pixelout<=1'b1;
2900: pixelout<=1'b1;
2901: pixelout<=1'b1;
2902: pixelout<=1'b1;
2903: pixelout<=1'b1;
2904: pixelout<=1'b1;
2905: pixelout<=1'b1;
2906: pixelout<=1'b1;
2907: pixelout<=1'b1;
2908: pixelout<=1'b1;
2909: pixelout<=1'b1;
2910: pixelout<=1'b1;
2911: pixelout<=1'b1;
2912: pixelout<=1'b1;
2913: pixelout<=1'b1;
2914: pixelout<=1'b1;
2915: pixelout<=1'b1;
2916: pixelout<=1'b1;
2917: pixelout<=1'b1;
2918: pixelout<=1'b1;
2919: pixelout<=1'b1;
2920: pixelout<=1'b1;
2921: pixelout<=1'b1;
2922: pixelout<=1'b1;
2923: pixelout<=1'b1;
2924: pixelout<=1'b1;
2925: pixelout<=1'b1;
2926: pixelout<=1'b1;
2927: pixelout<=1'b1;
2928: pixelout<=1'b1;
2929: pixelout<=1'b1;
2930: pixelout<=1'b0;
2931: pixelout<=1'b1;
2932: pixelout<=1'b1;
2933: pixelout<=1'b0;
2934: pixelout<=1'b0;
2935: pixelout<=1'b1;
2936: pixelout<=1'b1;
2937: pixelout<=1'b1;
2938: pixelout<=1'b1;
2939: pixelout<=1'b1;
2940: pixelout<=1'b1;
2941: pixelout<=1'b1;
2942: pixelout<=1'b1;
2943: pixelout<=1'b1;
2944: pixelout<=1'b1;
2945: pixelout<=1'b1;
2946: pixelout<=1'b1;
2947: pixelout<=1'b1;
2948: pixelout<=1'b1;
2949: pixelout<=1'b1;
2950: pixelout<=1'b1;
2951: pixelout<=1'b1;
2952: pixelout<=1'b1;
2953: pixelout<=1'b1;
2954: pixelout<=1'b1;
2955: pixelout<=1'b1;
2956: pixelout<=1'b1;
2957: pixelout<=1'b1;
2958: pixelout<=1'b1;
2959: pixelout<=1'b1;
2960: pixelout<=1'b1;
2961: pixelout<=1'b1;
2962: pixelout<=1'b1;
2963: pixelout<=1'b1;
2964: pixelout<=1'b1;
2965: pixelout<=1'b1;
2966: pixelout<=1'b1;
2967: pixelout<=1'b1;
2968: pixelout<=1'b1;
2969: pixelout<=1'b1;
2970: pixelout<=1'b1;
2971: pixelout<=1'b1;
2972: pixelout<=1'b1;
2973: pixelout<=1'b1;
2974: pixelout<=1'b1;
2975: pixelout<=1'b1;
2976: pixelout<=1'b1;
2977: pixelout<=1'b1;
2978: pixelout<=1'b1;
2979: pixelout<=1'b1;
2980: pixelout<=1'b1;
2981: pixelout<=1'b1;
2982: pixelout<=1'b0;
2983: pixelout<=1'b1;
2984: pixelout<=1'b1;
2985: pixelout<=1'b1;
2986: pixelout<=1'b1;
2987: pixelout<=1'b1;
2988: pixelout<=1'b1;
2989: pixelout<=1'b1;
2990: pixelout<=1'b1;
2991: pixelout<=1'b1;
2992: pixelout<=1'b1;
2993: pixelout<=1'b1;
2994: pixelout<=1'b1;
2995: pixelout<=1'b1;
2996: pixelout<=1'b1;
2997: pixelout<=1'b1;
2998: pixelout<=1'b1;
2999: pixelout<=1'b1;
3000: pixelout<=1'b1;
3001: pixelout<=1'b1;
3002: pixelout<=1'b1;
3003: pixelout<=1'b1;
3004: pixelout<=1'b1;
3005: pixelout<=1'b1;
3006: pixelout<=1'b1;
3007: pixelout<=1'b1;
3008: pixelout<=1'b1;
3009: pixelout<=1'b1;
3010: pixelout<=1'b1;
3011: pixelout<=1'b1;
3012: pixelout<=1'b1;
3013: pixelout<=1'b1;
3014: pixelout<=1'b1;
3015: pixelout<=1'b1;
3016: pixelout<=1'b1;
3017: pixelout<=1'b1;
3018: pixelout<=1'b1;
3019: pixelout<=1'b1;
3020: pixelout<=1'b1;
3021: pixelout<=1'b1;
3022: pixelout<=1'b1;
3023: pixelout<=1'b1;
3024: pixelout<=1'b1;
3025: pixelout<=1'b1;
3026: pixelout<=1'b1;
3027: pixelout<=1'b1;
3028: pixelout<=1'b1;
3029: pixelout<=1'b1;
3030: pixelout<=1'b1;
3031: pixelout<=1'b1;
3032: pixelout<=1'b1;
3033: pixelout<=1'b1;
3034: pixelout<=1'b1;
3035: pixelout<=1'b1;
3036: pixelout<=1'b1;
3037: pixelout<=1'b1;
3038: pixelout<=1'b1;
3039: pixelout<=1'b1;
3040: pixelout<=1'b1;
3041: pixelout<=1'b1;
3042: pixelout<=1'b1;
3043: pixelout<=1'b1;
3044: pixelout<=1'b1;
3045: pixelout<=1'b1;
3046: pixelout<=1'b1;
3047: pixelout<=1'b1;
3048: pixelout<=1'b1;
3049: pixelout<=1'b1;
3050: pixelout<=1'b1;
3051: pixelout<=1'b1;
3052: pixelout<=1'b1;
3053: pixelout<=1'b1;
3054: pixelout<=1'b1;
3055: pixelout<=1'b1;
3056: pixelout<=1'b1;
3057: pixelout<=1'b1;
3058: pixelout<=1'b1;
3059: pixelout<=1'b1;
3060: pixelout<=1'b1;
3061: pixelout<=1'b1;
3062: pixelout<=1'b1;
3063: pixelout<=1'b1;
3064: pixelout<=1'b1;
3065: pixelout<=1'b1;
3066: pixelout<=1'b1;
3067: pixelout<=1'b1;
3068: pixelout<=1'b1;
3069: pixelout<=1'b1;
3070: pixelout<=1'b1;
3071: pixelout<=1'b1;
3072: pixelout<=1'b1;
3073: pixelout<=1'b1;
3074: pixelout<=1'b1;
3075: pixelout<=1'b1;
3076: pixelout<=1'b1;
3077: pixelout<=1'b1;
3078: pixelout<=1'b1;
3079: pixelout<=1'b1;
3080: pixelout<=1'b1;
3081: pixelout<=1'b1;
3082: pixelout<=1'b1;
3083: pixelout<=1'b1;
3084: pixelout<=1'b1;
3085: pixelout<=1'b1;
3086: pixelout<=1'b0;
3087: pixelout<=1'b0;
3088: pixelout<=1'b0;
3089: pixelout<=1'b1;
3090: pixelout<=1'b1;
3091: pixelout<=1'b1;
3092: pixelout<=1'b1;
3093: pixelout<=1'b0;
3094: pixelout<=1'b0;
3095: pixelout<=1'b1;
3096: pixelout<=1'b1;
3097: pixelout<=1'b1;
3098: pixelout<=1'b0;
3099: pixelout<=1'b0;
3100: pixelout<=1'b0;
3101: pixelout<=1'b0;
3102: pixelout<=1'b1;
3103: pixelout<=1'b1;
3104: pixelout<=1'b1;
3105: pixelout<=1'b1;
3106: pixelout<=1'b1;
3107: pixelout<=1'b1;
3108: pixelout<=1'b1;
3109: pixelout<=1'b1;
3110: pixelout<=1'b1;
3111: pixelout<=1'b1;
3112: pixelout<=1'b1;
3113: pixelout<=1'b1;
3114: pixelout<=1'b1;
3115: pixelout<=1'b1;
3116: pixelout<=1'b1;
3117: pixelout<=1'b1;
3118: pixelout<=1'b1;
3119: pixelout<=1'b1;
3120: pixelout<=1'b1;
3121: pixelout<=1'b1;
3122: pixelout<=1'b1;
3123: pixelout<=1'b1;
3124: pixelout<=1'b1;
3125: pixelout<=1'b1;
3126: pixelout<=1'b1;
3127: pixelout<=1'b1;
3128: pixelout<=1'b1;
3129: pixelout<=1'b1;
3130: pixelout<=1'b1;
3131: pixelout<=1'b1;
3132: pixelout<=1'b1;
3133: pixelout<=1'b1;
3134: pixelout<=1'b1;
3135: pixelout<=1'b0;
3136: pixelout<=1'b0;
3137: pixelout<=1'b0;
3138: pixelout<=1'b0;
3139: pixelout<=1'b1;
3140: pixelout<=1'b1;
3141: pixelout<=1'b1;
3142: pixelout<=1'b1;
3143: pixelout<=1'b1;
3144: pixelout<=1'b1;
3145: pixelout<=1'b1;
3146: pixelout<=1'b1;
3147: pixelout<=1'b1;
3148: pixelout<=1'b1;
3149: pixelout<=1'b1;
3150: pixelout<=1'b1;
3151: pixelout<=1'b1;
3152: pixelout<=1'b1;
3153: pixelout<=1'b1;
3154: pixelout<=1'b1;
3155: pixelout<=1'b0;
3156: pixelout<=1'b0;
3157: pixelout<=1'b1;
3158: pixelout<=1'b1;
3159: pixelout<=1'b1;
3160: pixelout<=1'b1;
3161: pixelout<=1'b1;
3162: pixelout<=1'b1;
3163: pixelout<=1'b1;
3164: pixelout<=1'b1;
3165: pixelout<=1'b1;
3166: pixelout<=1'b1;
3167: pixelout<=1'b1;
3168: pixelout<=1'b1;
3169: pixelout<=1'b1;
3170: pixelout<=1'b1;
3171: pixelout<=1'b1;
3172: pixelout<=1'b1;
3173: pixelout<=1'b1;
3174: pixelout<=1'b1;
3175: pixelout<=1'b1;
3176: pixelout<=1'b1;
3177: pixelout<=1'b0;
3178: pixelout<=1'b0;
3179: pixelout<=1'b0;
3180: pixelout<=1'b1;
3181: pixelout<=1'b1;
3182: pixelout<=1'b1;
3183: pixelout<=1'b1;
3184: pixelout<=1'b1;
3185: pixelout<=1'b1;
3186: pixelout<=1'b1;
3187: pixelout<=1'b1;
3188: pixelout<=1'b1;
3189: pixelout<=1'b1;
3190: pixelout<=1'b1;
3191: pixelout<=1'b1;
3192: pixelout<=1'b1;
3193: pixelout<=1'b1;
3194: pixelout<=1'b1;
3195: pixelout<=1'b1;
3196: pixelout<=1'b1;
3197: pixelout<=1'b1;
3198: pixelout<=1'b1;
3199: pixelout<=1'b1;
3200: pixelout<=1'b1;
3201: pixelout<=1'b1;
3202: pixelout<=1'b1;
3203: pixelout<=1'b1;
3204: pixelout<=1'b1;
3205: pixelout<=1'b1;
3206: pixelout<=1'b1;
3207: pixelout<=1'b1;
3208: pixelout<=1'b1;
3209: pixelout<=1'b1;
3210: pixelout<=1'b1;
3211: pixelout<=1'b1;
3212: pixelout<=1'b1;
3213: pixelout<=1'b1;
3214: pixelout<=1'b1;
3215: pixelout<=1'b1;
3216: pixelout<=1'b1;
3217: pixelout<=1'b1;
3218: pixelout<=1'b1;
3219: pixelout<=1'b1;
3220: pixelout<=1'b1;
3221: pixelout<=1'b1;
3222: pixelout<=1'b0;
3223: pixelout<=1'b1;
3224: pixelout<=1'b1;
3225: pixelout<=1'b1;
3226: pixelout<=1'b0;
3227: pixelout<=1'b1;
3228: pixelout<=1'b1;
3229: pixelout<=1'b1;
3230: pixelout<=1'b0;
3231: pixelout<=1'b1;
3232: pixelout<=1'b1;
3233: pixelout<=1'b1;
3234: pixelout<=1'b1;
3235: pixelout<=1'b1;
3236: pixelout<=1'b1;
3237: pixelout<=1'b1;
3238: pixelout<=1'b1;
3239: pixelout<=1'b1;
3240: pixelout<=1'b1;
3241: pixelout<=1'b1;
3242: pixelout<=1'b1;
3243: pixelout<=1'b1;
3244: pixelout<=1'b1;
3245: pixelout<=1'b1;
3246: pixelout<=1'b1;
3247: pixelout<=1'b1;
3248: pixelout<=1'b1;
3249: pixelout<=1'b1;
3250: pixelout<=1'b1;
3251: pixelout<=1'b1;
3252: pixelout<=1'b1;
3253: pixelout<=1'b1;
3254: pixelout<=1'b1;
3255: pixelout<=1'b1;
3256: pixelout<=1'b1;
3257: pixelout<=1'b1;
3258: pixelout<=1'b1;
3259: pixelout<=1'b1;
3260: pixelout<=1'b1;
3261: pixelout<=1'b1;
3262: pixelout<=1'b1;
3263: pixelout<=1'b1;
3264: pixelout<=1'b1;
3265: pixelout<=1'b1;
3266: pixelout<=1'b1;
3267: pixelout<=1'b1;
3268: pixelout<=1'b1;
3269: pixelout<=1'b1;
3270: pixelout<=1'b1;
3271: pixelout<=1'b1;
3272: pixelout<=1'b1;
3273: pixelout<=1'b1;
3274: pixelout<=1'b1;
3275: pixelout<=1'b1;
3276: pixelout<=1'b1;
3277: pixelout<=1'b1;
3278: pixelout<=1'b1;
3279: pixelout<=1'b1;
3280: pixelout<=1'b1;
3281: pixelout<=1'b1;
3282: pixelout<=1'b0;
3283: pixelout<=1'b0;
3284: pixelout<=1'b1;
3285: pixelout<=1'b1;
3286: pixelout<=1'b1;
3287: pixelout<=1'b1;
3288: pixelout<=1'b1;
3289: pixelout<=1'b1;
3290: pixelout<=1'b1;
3291: pixelout<=1'b1;
3292: pixelout<=1'b1;
3293: pixelout<=1'b1;
3294: pixelout<=1'b1;
3295: pixelout<=1'b1;
3296: pixelout<=1'b1;
3297: pixelout<=1'b1;
3298: pixelout<=1'b1;
3299: pixelout<=1'b1;
3300: pixelout<=1'b1;
3301: pixelout<=1'b1;
3302: pixelout<=1'b1;
3303: pixelout<=1'b1;
3304: pixelout<=1'b0;
3305: pixelout<=1'b0;
3306: pixelout<=1'b0;
3307: pixelout<=1'b0;
3308: pixelout<=1'b0;
3309: pixelout<=1'b1;
3310: pixelout<=1'b1;
3311: pixelout<=1'b1;
3312: pixelout<=1'b0;
3313: pixelout<=1'b0;
3314: pixelout<=1'b1;
3315: pixelout<=1'b1;
3316: pixelout<=1'b1;
3317: pixelout<=1'b0;
3318: pixelout<=1'b0;
3319: pixelout<=1'b0;
3320: pixelout<=1'b0;
3321: pixelout<=1'b1;
3322: pixelout<=1'b1;
3323: pixelout<=1'b1;
3324: pixelout<=1'b1;
3325: pixelout<=1'b0;
3326: pixelout<=1'b1;
3327: pixelout<=1'b1;
3328: pixelout<=1'b1;
3329: pixelout<=1'b0;
3330: pixelout<=1'b1;
3331: pixelout<=1'b0;
3332: pixelout<=1'b1;
3333: pixelout<=1'b1;
3334: pixelout<=1'b1;
3335: pixelout<=1'b1;
3336: pixelout<=1'b1;
3337: pixelout<=1'b1;
3338: pixelout<=1'b1;
3339: pixelout<=1'b1;
3340: pixelout<=1'b1;
3341: pixelout<=1'b1;
3342: pixelout<=1'b1;
3343: pixelout<=1'b1;
3344: pixelout<=1'b1;
3345: pixelout<=1'b1;
3346: pixelout<=1'b1;
3347: pixelout<=1'b1;
3348: pixelout<=1'b1;
3349: pixelout<=1'b1;
3350: pixelout<=1'b1;
3351: pixelout<=1'b1;
3352: pixelout<=1'b1;
3353: pixelout<=1'b1;
3354: pixelout<=1'b1;
3355: pixelout<=1'b1;
3356: pixelout<=1'b1;
3357: pixelout<=1'b1;
3358: pixelout<=1'b1;
3359: pixelout<=1'b1;
3360: pixelout<=1'b1;
3361: pixelout<=1'b1;
3362: pixelout<=1'b1;
3363: pixelout<=1'b1;
3364: pixelout<=1'b1;
3365: pixelout<=1'b1;
3366: pixelout<=1'b1;
3367: pixelout<=1'b1;
3368: pixelout<=1'b1;
3369: pixelout<=1'b1;
3370: pixelout<=1'b1;
3371: pixelout<=1'b1;
3372: pixelout<=1'b1;
3373: pixelout<=1'b1;
3374: pixelout<=1'b1;
3375: pixelout<=1'b1;
3376: pixelout<=1'b1;
3377: pixelout<=1'b1;
3378: pixelout<=1'b1;
3379: pixelout<=1'b1;
3380: pixelout<=1'b1;
3381: pixelout<=1'b1;
3382: pixelout<=1'b1;
3383: pixelout<=1'b1;
3384: pixelout<=1'b1;
3385: pixelout<=1'b1;
3386: pixelout<=1'b1;
3387: pixelout<=1'b1;
3388: pixelout<=1'b1;
3389: pixelout<=1'b1;
3390: pixelout<=1'b1;
3391: pixelout<=1'b1;
3392: pixelout<=1'b1;
3393: pixelout<=1'b1;
3394: pixelout<=1'b0;
3395: pixelout<=1'b1;
3396: pixelout<=1'b1;
3397: pixelout<=1'b1;
3398: pixelout<=1'b1;
3399: pixelout<=1'b1;
3400: pixelout<=1'b1;
3401: pixelout<=1'b1;
3402: pixelout<=1'b1;
3403: pixelout<=1'b1;
3404: pixelout<=1'b1;
3405: pixelout<=1'b0;
3406: pixelout<=1'b1;
3407: pixelout<=1'b1;
3408: pixelout<=1'b1;
3409: pixelout<=1'b1;
3410: pixelout<=1'b1;
3411: pixelout<=1'b1;
3412: pixelout<=1'b1;
3413: pixelout<=1'b1;
3414: pixelout<=1'b1;
3415: pixelout<=1'b1;
3416: pixelout<=1'b0;
3417: pixelout<=1'b1;
3418: pixelout<=1'b1;
3419: pixelout<=1'b1;
3420: pixelout<=1'b1;
3421: pixelout<=1'b1;
3422: pixelout<=1'b1;
3423: pixelout<=1'b1;
3424: pixelout<=1'b1;
3425: pixelout<=1'b1;
3426: pixelout<=1'b1;
3427: pixelout<=1'b1;
3428: pixelout<=1'b1;
3429: pixelout<=1'b1;
3430: pixelout<=1'b1;
3431: pixelout<=1'b1;
3432: pixelout<=1'b1;
3433: pixelout<=1'b1;
3434: pixelout<=1'b1;
3435: pixelout<=1'b1;
3436: pixelout<=1'b1;
3437: pixelout<=1'b1;
3438: pixelout<=1'b1;
3439: pixelout<=1'b1;
3440: pixelout<=1'b1;
3441: pixelout<=1'b1;
3442: pixelout<=1'b1;
3443: pixelout<=1'b1;
3444: pixelout<=1'b1;
3445: pixelout<=1'b1;
3446: pixelout<=1'b1;
3447: pixelout<=1'b1;
3448: pixelout<=1'b1;
3449: pixelout<=1'b1;
3450: pixelout<=1'b1;
3451: pixelout<=1'b1;
3452: pixelout<=1'b1;
3453: pixelout<=1'b1;
3454: pixelout<=1'b1;
3455: pixelout<=1'b1;
3456: pixelout<=1'b1;
3457: pixelout<=1'b1;
3458: pixelout<=1'b1;
3459: pixelout<=1'b1;
3460: pixelout<=1'b1;
3461: pixelout<=1'b1;
3462: pixelout<=1'b0;
3463: pixelout<=1'b1;
3464: pixelout<=1'b1;
3465: pixelout<=1'b1;
3466: pixelout<=1'b0;
3467: pixelout<=1'b1;
3468: pixelout<=1'b1;
3469: pixelout<=1'b1;
3470: pixelout<=1'b1;
3471: pixelout<=1'b1;
3472: pixelout<=1'b1;
3473: pixelout<=1'b1;
3474: pixelout<=1'b1;
3475: pixelout<=1'b1;
3476: pixelout<=1'b1;
3477: pixelout<=1'b1;
3478: pixelout<=1'b1;
3479: pixelout<=1'b1;
3480: pixelout<=1'b1;
3481: pixelout<=1'b1;
3482: pixelout<=1'b1;
3483: pixelout<=1'b1;
3484: pixelout<=1'b1;
3485: pixelout<=1'b1;
3486: pixelout<=1'b1;
3487: pixelout<=1'b1;
3488: pixelout<=1'b1;
3489: pixelout<=1'b1;
3490: pixelout<=1'b1;
3491: pixelout<=1'b1;
3492: pixelout<=1'b1;
3493: pixelout<=1'b1;
3494: pixelout<=1'b1;
3495: pixelout<=1'b1;
3496: pixelout<=1'b1;
3497: pixelout<=1'b1;
3498: pixelout<=1'b1;
3499: pixelout<=1'b1;
3500: pixelout<=1'b0;
3501: pixelout<=1'b1;
3502: pixelout<=1'b1;
3503: pixelout<=1'b1;
3504: pixelout<=1'b1;
3505: pixelout<=1'b1;
3506: pixelout<=1'b1;
3507: pixelout<=1'b1;
3508: pixelout<=1'b1;
3509: pixelout<=1'b1;
3510: pixelout<=1'b1;
3511: pixelout<=1'b1;
3512: pixelout<=1'b1;
3513: pixelout<=1'b1;
3514: pixelout<=1'b1;
3515: pixelout<=1'b1;
3516: pixelout<=1'b1;
3517: pixelout<=1'b1;
3518: pixelout<=1'b1;
3519: pixelout<=1'b1;
3520: pixelout<=1'b0;
3521: pixelout<=1'b1;
3522: pixelout<=1'b1;
3523: pixelout<=1'b1;
3524: pixelout<=1'b1;
3525: pixelout<=1'b1;
3526: pixelout<=1'b1;
3527: pixelout<=1'b1;
3528: pixelout<=1'b1;
3529: pixelout<=1'b0;
3530: pixelout<=1'b1;
3531: pixelout<=1'b1;
3532: pixelout<=1'b1;
3533: pixelout<=1'b1;
3534: pixelout<=1'b1;
3535: pixelout<=1'b1;
3536: pixelout<=1'b1;
3537: pixelout<=1'b1;
3538: pixelout<=1'b1;
3539: pixelout<=1'b1;
3540: pixelout<=1'b1;
3541: pixelout<=1'b1;
3542: pixelout<=1'b1;
3543: pixelout<=1'b1;
3544: pixelout<=1'b0;
3545: pixelout<=1'b1;
3546: pixelout<=1'b1;
3547: pixelout<=1'b1;
3548: pixelout<=1'b1;
3549: pixelout<=1'b1;
3550: pixelout<=1'b0;
3551: pixelout<=1'b1;
3552: pixelout<=1'b1;
3553: pixelout<=1'b1;
3554: pixelout<=1'b1;
3555: pixelout<=1'b1;
3556: pixelout<=1'b1;
3557: pixelout<=1'b1;
3558: pixelout<=1'b1;
3559: pixelout<=1'b1;
3560: pixelout<=1'b1;
3561: pixelout<=1'b1;
3562: pixelout<=1'b1;
3563: pixelout<=1'b1;
3564: pixelout<=1'b1;
3565: pixelout<=1'b1;
3566: pixelout<=1'b1;
3567: pixelout<=1'b1;
3568: pixelout<=1'b1;
3569: pixelout<=1'b0;
3570: pixelout<=1'b1;
3571: pixelout<=1'b0;
3572: pixelout<=1'b1;
3573: pixelout<=1'b1;
3574: pixelout<=1'b1;
3575: pixelout<=1'b1;
3576: pixelout<=1'b1;
3577: pixelout<=1'b1;
3578: pixelout<=1'b1;
3579: pixelout<=1'b1;
3580: pixelout<=1'b1;
3581: pixelout<=1'b1;
3582: pixelout<=1'b1;
3583: pixelout<=1'b1;
3584: pixelout<=1'b1;
3585: pixelout<=1'b1;
3586: pixelout<=1'b1;
3587: pixelout<=1'b1;
3588: pixelout<=1'b1;
3589: pixelout<=1'b1;
3590: pixelout<=1'b1;
3591: pixelout<=1'b1;
3592: pixelout<=1'b1;
3593: pixelout<=1'b1;
3594: pixelout<=1'b1;
3595: pixelout<=1'b1;
3596: pixelout<=1'b1;
3597: pixelout<=1'b1;
3598: pixelout<=1'b1;
3599: pixelout<=1'b1;
3600: pixelout<=1'b1;
3601: pixelout<=1'b1;
3602: pixelout<=1'b1;
3603: pixelout<=1'b1;
3604: pixelout<=1'b1;
3605: pixelout<=1'b1;
3606: pixelout<=1'b1;
3607: pixelout<=1'b1;
3608: pixelout<=1'b1;
3609: pixelout<=1'b1;
3610: pixelout<=1'b1;
3611: pixelout<=1'b1;
3612: pixelout<=1'b1;
3613: pixelout<=1'b1;
3614: pixelout<=1'b1;
3615: pixelout<=1'b1;
3616: pixelout<=1'b1;
3617: pixelout<=1'b1;
3618: pixelout<=1'b1;
3619: pixelout<=1'b1;
3620: pixelout<=1'b1;
3621: pixelout<=1'b1;
3622: pixelout<=1'b1;
3623: pixelout<=1'b1;
3624: pixelout<=1'b1;
3625: pixelout<=1'b1;
3626: pixelout<=1'b1;
3627: pixelout<=1'b1;
3628: pixelout<=1'b1;
3629: pixelout<=1'b1;
3630: pixelout<=1'b1;
3631: pixelout<=1'b1;
3632: pixelout<=1'b1;
3633: pixelout<=1'b1;
3634: pixelout<=1'b0;
3635: pixelout<=1'b1;
3636: pixelout<=1'b1;
3637: pixelout<=1'b1;
3638: pixelout<=1'b1;
3639: pixelout<=1'b1;
3640: pixelout<=1'b1;
3641: pixelout<=1'b1;
3642: pixelout<=1'b1;
3643: pixelout<=1'b1;
3644: pixelout<=1'b1;
3645: pixelout<=1'b0;
3646: pixelout<=1'b1;
3647: pixelout<=1'b1;
3648: pixelout<=1'b1;
3649: pixelout<=1'b1;
3650: pixelout<=1'b1;
3651: pixelout<=1'b1;
3652: pixelout<=1'b1;
3653: pixelout<=1'b1;
3654: pixelout<=1'b1;
3655: pixelout<=1'b1;
3656: pixelout<=1'b0;
3657: pixelout<=1'b1;
3658: pixelout<=1'b1;
3659: pixelout<=1'b1;
3660: pixelout<=1'b1;
3661: pixelout<=1'b1;
3662: pixelout<=1'b1;
3663: pixelout<=1'b1;
3664: pixelout<=1'b1;
3665: pixelout<=1'b1;
3666: pixelout<=1'b1;
3667: pixelout<=1'b1;
3668: pixelout<=1'b1;
3669: pixelout<=1'b1;
3670: pixelout<=1'b1;
3671: pixelout<=1'b1;
3672: pixelout<=1'b1;
3673: pixelout<=1'b1;
3674: pixelout<=1'b1;
3675: pixelout<=1'b1;
3676: pixelout<=1'b1;
3677: pixelout<=1'b1;
3678: pixelout<=1'b1;
3679: pixelout<=1'b1;
3680: pixelout<=1'b1;
3681: pixelout<=1'b1;
3682: pixelout<=1'b1;
3683: pixelout<=1'b1;
3684: pixelout<=1'b1;
3685: pixelout<=1'b1;
3686: pixelout<=1'b1;
3687: pixelout<=1'b1;
3688: pixelout<=1'b1;
3689: pixelout<=1'b1;
3690: pixelout<=1'b1;
3691: pixelout<=1'b1;
3692: pixelout<=1'b1;
3693: pixelout<=1'b1;
3694: pixelout<=1'b1;
3695: pixelout<=1'b1;
3696: pixelout<=1'b1;
3697: pixelout<=1'b1;
3698: pixelout<=1'b1;
3699: pixelout<=1'b1;
3700: pixelout<=1'b1;
3701: pixelout<=1'b1;
3702: pixelout<=1'b0;
3703: pixelout<=1'b1;
3704: pixelout<=1'b1;
3705: pixelout<=1'b1;
3706: pixelout<=1'b1;
3707: pixelout<=1'b0;
3708: pixelout<=1'b1;
3709: pixelout<=1'b0;
3710: pixelout<=1'b1;
3711: pixelout<=1'b1;
3712: pixelout<=1'b1;
3713: pixelout<=1'b1;
3714: pixelout<=1'b1;
3715: pixelout<=1'b1;
3716: pixelout<=1'b1;
3717: pixelout<=1'b1;
3718: pixelout<=1'b1;
3719: pixelout<=1'b1;
3720: pixelout<=1'b1;
3721: pixelout<=1'b1;
3722: pixelout<=1'b1;
3723: pixelout<=1'b1;
3724: pixelout<=1'b1;
3725: pixelout<=1'b1;
3726: pixelout<=1'b1;
3727: pixelout<=1'b1;
3728: pixelout<=1'b1;
3729: pixelout<=1'b1;
3730: pixelout<=1'b1;
3731: pixelout<=1'b1;
3732: pixelout<=1'b1;
3733: pixelout<=1'b1;
3734: pixelout<=1'b1;
3735: pixelout<=1'b1;
3736: pixelout<=1'b1;
3737: pixelout<=1'b1;
3738: pixelout<=1'b1;
3739: pixelout<=1'b1;
3740: pixelout<=1'b0;
3741: pixelout<=1'b1;
3742: pixelout<=1'b1;
3743: pixelout<=1'b1;
3744: pixelout<=1'b1;
3745: pixelout<=1'b1;
3746: pixelout<=1'b1;
3747: pixelout<=1'b1;
3748: pixelout<=1'b1;
3749: pixelout<=1'b1;
3750: pixelout<=1'b1;
3751: pixelout<=1'b1;
3752: pixelout<=1'b1;
3753: pixelout<=1'b1;
3754: pixelout<=1'b1;
3755: pixelout<=1'b1;
3756: pixelout<=1'b1;
3757: pixelout<=1'b1;
3758: pixelout<=1'b1;
3759: pixelout<=1'b1;
3760: pixelout<=1'b0;
3761: pixelout<=1'b1;
3762: pixelout<=1'b1;
3763: pixelout<=1'b1;
3764: pixelout<=1'b1;
3765: pixelout<=1'b1;
3766: pixelout<=1'b1;
3767: pixelout<=1'b1;
3768: pixelout<=1'b1;
3769: pixelout<=1'b0;
3770: pixelout<=1'b1;
3771: pixelout<=1'b1;
3772: pixelout<=1'b1;
3773: pixelout<=1'b1;
3774: pixelout<=1'b1;
3775: pixelout<=1'b1;
3776: pixelout<=1'b1;
3777: pixelout<=1'b1;
3778: pixelout<=1'b1;
3779: pixelout<=1'b1;
3780: pixelout<=1'b1;
3781: pixelout<=1'b1;
3782: pixelout<=1'b1;
3783: pixelout<=1'b1;
3784: pixelout<=1'b0;
3785: pixelout<=1'b1;
3786: pixelout<=1'b1;
3787: pixelout<=1'b1;
3788: pixelout<=1'b1;
3789: pixelout<=1'b1;
3790: pixelout<=1'b0;
3791: pixelout<=1'b1;
3792: pixelout<=1'b1;
3793: pixelout<=1'b1;
3794: pixelout<=1'b1;
3795: pixelout<=1'b1;
3796: pixelout<=1'b1;
3797: pixelout<=1'b1;
3798: pixelout<=1'b1;
3799: pixelout<=1'b1;
3800: pixelout<=1'b1;
3801: pixelout<=1'b1;
3802: pixelout<=1'b1;
3803: pixelout<=1'b1;
3804: pixelout<=1'b1;
3805: pixelout<=1'b1;
3806: pixelout<=1'b1;
3807: pixelout<=1'b1;
3808: pixelout<=1'b1;
3809: pixelout<=1'b1;
3810: pixelout<=1'b1;
3811: pixelout<=1'b1;
3812: pixelout<=1'b1;
3813: pixelout<=1'b1;
3814: pixelout<=1'b1;
3815: pixelout<=1'b1;
3816: pixelout<=1'b1;
3817: pixelout<=1'b1;
3818: pixelout<=1'b1;
3819: pixelout<=1'b1;
3820: pixelout<=1'b1;
3821: pixelout<=1'b1;
3822: pixelout<=1'b1;
3823: pixelout<=1'b1;
3824: pixelout<=1'b1;
3825: pixelout<=1'b1;
3826: pixelout<=1'b1;
3827: pixelout<=1'b1;
3828: pixelout<=1'b1;
3829: pixelout<=1'b1;
3830: pixelout<=1'b1;
3831: pixelout<=1'b1;
3832: pixelout<=1'b1;
3833: pixelout<=1'b1;
3834: pixelout<=1'b1;
3835: pixelout<=1'b1;
3836: pixelout<=1'b1;
3837: pixelout<=1'b1;
3838: pixelout<=1'b1;
3839: pixelout<=1'b1;
3840: pixelout<=1'b1;
3841: pixelout<=1'b1;
3842: pixelout<=1'b1;
3843: pixelout<=1'b1;
3844: pixelout<=1'b1;
3845: pixelout<=1'b1;
3846: pixelout<=1'b1;
3847: pixelout<=1'b1;
3848: pixelout<=1'b1;
3849: pixelout<=1'b1;
3850: pixelout<=1'b1;
3851: pixelout<=1'b1;
3852: pixelout<=1'b1;
3853: pixelout<=1'b1;
3854: pixelout<=1'b1;
3855: pixelout<=1'b1;
3856: pixelout<=1'b0;
3857: pixelout<=1'b1;
3858: pixelout<=1'b1;
3859: pixelout<=1'b1;
3860: pixelout<=1'b1;
3861: pixelout<=1'b1;
3862: pixelout<=1'b1;
3863: pixelout<=1'b1;
3864: pixelout<=1'b0;
3865: pixelout<=1'b1;
3866: pixelout<=1'b1;
3867: pixelout<=1'b1;
3868: pixelout<=1'b0;
3869: pixelout<=1'b0;
3870: pixelout<=1'b0;
3871: pixelout<=1'b1;
3872: pixelout<=1'b1;
3873: pixelout<=1'b0;
3874: pixelout<=1'b0;
3875: pixelout<=1'b0;
3876: pixelout<=1'b0;
3877: pixelout<=1'b1;
3878: pixelout<=1'b0;
3879: pixelout<=1'b1;
3880: pixelout<=1'b1;
3881: pixelout<=1'b0;
3882: pixelout<=1'b1;
3883: pixelout<=1'b1;
3884: pixelout<=1'b1;
3885: pixelout<=1'b1;
3886: pixelout<=1'b1;
3887: pixelout<=1'b1;
3888: pixelout<=1'b1;
3889: pixelout<=1'b1;
3890: pixelout<=1'b1;
3891: pixelout<=1'b1;
3892: pixelout<=1'b1;
3893: pixelout<=1'b1;
3894: pixelout<=1'b1;
3895: pixelout<=1'b1;
3896: pixelout<=1'b0;
3897: pixelout<=1'b1;
3898: pixelout<=1'b1;
3899: pixelout<=1'b1;
3900: pixelout<=1'b1;
3901: pixelout<=1'b1;
3902: pixelout<=1'b1;
3903: pixelout<=1'b1;
3904: pixelout<=1'b0;
3905: pixelout<=1'b0;
3906: pixelout<=1'b1;
3907: pixelout<=1'b1;
3908: pixelout<=1'b1;
3909: pixelout<=1'b0;
3910: pixelout<=1'b0;
3911: pixelout<=1'b1;
3912: pixelout<=1'b1;
3913: pixelout<=1'b1;
3914: pixelout<=1'b1;
3915: pixelout<=1'b0;
3916: pixelout<=1'b0;
3917: pixelout<=1'b0;
3918: pixelout<=1'b1;
3919: pixelout<=1'b1;
3920: pixelout<=1'b0;
3921: pixelout<=1'b1;
3922: pixelout<=1'b0;
3923: pixelout<=1'b0;
3924: pixelout<=1'b1;
3925: pixelout<=1'b1;
3926: pixelout<=1'b1;
3927: pixelout<=1'b0;
3928: pixelout<=1'b0;
3929: pixelout<=1'b0;
3930: pixelout<=1'b1;
3931: pixelout<=1'b1;
3932: pixelout<=1'b0;
3933: pixelout<=1'b0;
3934: pixelout<=1'b0;
3935: pixelout<=1'b1;
3936: pixelout<=1'b1;
3937: pixelout<=1'b0;
3938: pixelout<=1'b0;
3939: pixelout<=1'b0;
3940: pixelout<=1'b1;
3941: pixelout<=1'b1;
3942: pixelout<=1'b0;
3943: pixelout<=1'b1;
3944: pixelout<=1'b1;
3945: pixelout<=1'b1;
3946: pixelout<=1'b1;
3947: pixelout<=1'b0;
3948: pixelout<=1'b1;
3949: pixelout<=1'b0;
3950: pixelout<=1'b1;
3951: pixelout<=1'b1;
3952: pixelout<=1'b1;
3953: pixelout<=1'b1;
3954: pixelout<=1'b0;
3955: pixelout<=1'b0;
3956: pixelout<=1'b1;
3957: pixelout<=1'b1;
3958: pixelout<=1'b1;
3959: pixelout<=1'b1;
3960: pixelout<=1'b1;
3961: pixelout<=1'b1;
3962: pixelout<=1'b0;
3963: pixelout<=1'b1;
3964: pixelout<=1'b1;
3965: pixelout<=1'b1;
3966: pixelout<=1'b1;
3967: pixelout<=1'b1;
3968: pixelout<=1'b0;
3969: pixelout<=1'b0;
3970: pixelout<=1'b0;
3971: pixelout<=1'b1;
3972: pixelout<=1'b1;
3973: pixelout<=1'b1;
3974: pixelout<=1'b0;
3975: pixelout<=1'b0;
3976: pixelout<=1'b0;
3977: pixelout<=1'b1;
3978: pixelout<=1'b1;
3979: pixelout<=1'b1;
3980: pixelout<=1'b0;
3981: pixelout<=1'b0;
3982: pixelout<=1'b0;
3983: pixelout<=1'b1;
3984: pixelout<=1'b1;
3985: pixelout<=1'b1;
3986: pixelout<=1'b1;
3987: pixelout<=1'b1;
3988: pixelout<=1'b0;
3989: pixelout<=1'b0;
3990: pixelout<=1'b0;
3991: pixelout<=1'b0;
3992: pixelout<=1'b1;
3993: pixelout<=1'b0;
3994: pixelout<=1'b0;
3995: pixelout<=1'b0;
3996: pixelout<=1'b1;
3997: pixelout<=1'b1;
3998: pixelout<=1'b1;
3999: pixelout<=1'b1;
4000: pixelout<=1'b0;
4001: pixelout<=1'b1;
4002: pixelout<=1'b1;
4003: pixelout<=1'b1;
4004: pixelout<=1'b1;
4005: pixelout<=1'b1;
4006: pixelout<=1'b1;
4007: pixelout<=1'b0;
4008: pixelout<=1'b0;
4009: pixelout<=1'b0;
4010: pixelout<=1'b0;
4011: pixelout<=1'b1;
4012: pixelout<=1'b1;
4013: pixelout<=1'b1;
4014: pixelout<=1'b1;
4015: pixelout<=1'b0;
4016: pixelout<=1'b1;
4017: pixelout<=1'b0;
4018: pixelout<=1'b0;
4019: pixelout<=1'b0;
4020: pixelout<=1'b1;
4021: pixelout<=1'b1;
4022: pixelout<=1'b1;
4023: pixelout<=1'b1;
4024: pixelout<=1'b0;
4025: pixelout<=1'b0;
4026: pixelout<=1'b0;
4027: pixelout<=1'b0;
4028: pixelout<=1'b1;
4029: pixelout<=1'b1;
4030: pixelout<=1'b0;
4031: pixelout<=1'b1;
4032: pixelout<=1'b1;
4033: pixelout<=1'b1;
4034: pixelout<=1'b1;
4035: pixelout<=1'b1;
4036: pixelout<=1'b1;
4037: pixelout<=1'b0;
4038: pixelout<=1'b0;
4039: pixelout<=1'b0;
4040: pixelout<=1'b1;
4041: pixelout<=1'b1;
4042: pixelout<=1'b1;
4043: pixelout<=1'b1;
4044: pixelout<=1'b1;
4045: pixelout<=1'b1;
4046: pixelout<=1'b1;
4047: pixelout<=1'b0;
4048: pixelout<=1'b0;
4049: pixelout<=1'b1;
4050: pixelout<=1'b1;
4051: pixelout<=1'b1;
4052: pixelout<=1'b1;
4053: pixelout<=1'b0;
4054: pixelout<=1'b0;
4055: pixelout<=1'b1;
4056: pixelout<=1'b1;
4057: pixelout<=1'b1;
4058: pixelout<=1'b0;
4059: pixelout<=1'b0;
4060: pixelout<=1'b0;
4061: pixelout<=1'b1;
4062: pixelout<=1'b1;
4063: pixelout<=1'b1;
4064: pixelout<=1'b1;
4065: pixelout<=1'b1;
4066: pixelout<=1'b1;
4067: pixelout<=1'b1;
4068: pixelout<=1'b1;
4069: pixelout<=1'b1;
4070: pixelout<=1'b1;
4071: pixelout<=1'b1;
4072: pixelout<=1'b1;
4073: pixelout<=1'b1;
4074: pixelout<=1'b1;
4075: pixelout<=1'b1;
4076: pixelout<=1'b1;
4077: pixelout<=1'b1;
4078: pixelout<=1'b1;
4079: pixelout<=1'b1;
4080: pixelout<=1'b1;
4081: pixelout<=1'b1;
4082: pixelout<=1'b1;
4083: pixelout<=1'b1;
4084: pixelout<=1'b1;
4085: pixelout<=1'b1;
4086: pixelout<=1'b1;
4087: pixelout<=1'b1;
4088: pixelout<=1'b1;
4089: pixelout<=1'b1;
4090: pixelout<=1'b1;
4091: pixelout<=1'b1;
4092: pixelout<=1'b1;
4093: pixelout<=1'b1;
4094: pixelout<=1'b1;
4095: pixelout<=1'b1;
4096: pixelout<=1'b0;
4097: pixelout<=1'b1;
4098: pixelout<=1'b1;
4099: pixelout<=1'b1;
4100: pixelout<=1'b1;
4101: pixelout<=1'b1;
4102: pixelout<=1'b1;
4103: pixelout<=1'b1;
4104: pixelout<=1'b0;
4105: pixelout<=1'b1;
4106: pixelout<=1'b1;
4107: pixelout<=1'b0;
4108: pixelout<=1'b1;
4109: pixelout<=1'b1;
4110: pixelout<=1'b1;
4111: pixelout<=1'b0;
4112: pixelout<=1'b1;
4113: pixelout<=1'b1;
4114: pixelout<=1'b0;
4115: pixelout<=1'b1;
4116: pixelout<=1'b1;
4117: pixelout<=1'b1;
4118: pixelout<=1'b0;
4119: pixelout<=1'b1;
4120: pixelout<=1'b1;
4121: pixelout<=1'b0;
4122: pixelout<=1'b1;
4123: pixelout<=1'b1;
4124: pixelout<=1'b1;
4125: pixelout<=1'b1;
4126: pixelout<=1'b1;
4127: pixelout<=1'b1;
4128: pixelout<=1'b1;
4129: pixelout<=1'b1;
4130: pixelout<=1'b1;
4131: pixelout<=1'b1;
4132: pixelout<=1'b1;
4133: pixelout<=1'b1;
4134: pixelout<=1'b1;
4135: pixelout<=1'b1;
4136: pixelout<=1'b0;
4137: pixelout<=1'b1;
4138: pixelout<=1'b1;
4139: pixelout<=1'b1;
4140: pixelout<=1'b1;
4141: pixelout<=1'b1;
4142: pixelout<=1'b0;
4143: pixelout<=1'b1;
4144: pixelout<=1'b1;
4145: pixelout<=1'b1;
4146: pixelout<=1'b1;
4147: pixelout<=1'b1;
4148: pixelout<=1'b1;
4149: pixelout<=1'b1;
4150: pixelout<=1'b1;
4151: pixelout<=1'b1;
4152: pixelout<=1'b0;
4153: pixelout<=1'b1;
4154: pixelout<=1'b0;
4155: pixelout<=1'b1;
4156: pixelout<=1'b1;
4157: pixelout<=1'b1;
4158: pixelout<=1'b0;
4159: pixelout<=1'b1;
4160: pixelout<=1'b0;
4161: pixelout<=1'b0;
4162: pixelout<=1'b1;
4163: pixelout<=1'b1;
4164: pixelout<=1'b1;
4165: pixelout<=1'b0;
4166: pixelout<=1'b1;
4167: pixelout<=1'b1;
4168: pixelout<=1'b1;
4169: pixelout<=1'b1;
4170: pixelout<=1'b1;
4171: pixelout<=1'b1;
4172: pixelout<=1'b1;
4173: pixelout<=1'b1;
4174: pixelout<=1'b1;
4175: pixelout<=1'b1;
4176: pixelout<=1'b1;
4177: pixelout<=1'b1;
4178: pixelout<=1'b1;
4179: pixelout<=1'b1;
4180: pixelout<=1'b1;
4181: pixelout<=1'b1;
4182: pixelout<=1'b0;
4183: pixelout<=1'b1;
4184: pixelout<=1'b1;
4185: pixelout<=1'b1;
4186: pixelout<=1'b1;
4187: pixelout<=1'b1;
4188: pixelout<=1'b0;
4189: pixelout<=1'b1;
4190: pixelout<=1'b1;
4191: pixelout<=1'b1;
4192: pixelout<=1'b0;
4193: pixelout<=1'b1;
4194: pixelout<=1'b1;
4195: pixelout<=1'b1;
4196: pixelout<=1'b1;
4197: pixelout<=1'b1;
4198: pixelout<=1'b1;
4199: pixelout<=1'b1;
4200: pixelout<=1'b1;
4201: pixelout<=1'b1;
4202: pixelout<=1'b0;
4203: pixelout<=1'b1;
4204: pixelout<=1'b1;
4205: pixelout<=1'b1;
4206: pixelout<=1'b1;
4207: pixelout<=1'b0;
4208: pixelout<=1'b1;
4209: pixelout<=1'b1;
4210: pixelout<=1'b1;
4211: pixelout<=1'b0;
4212: pixelout<=1'b1;
4213: pixelout<=1'b0;
4214: pixelout<=1'b1;
4215: pixelout<=1'b1;
4216: pixelout<=1'b1;
4217: pixelout<=1'b0;
4218: pixelout<=1'b1;
4219: pixelout<=1'b1;
4220: pixelout<=1'b0;
4221: pixelout<=1'b1;
4222: pixelout<=1'b1;
4223: pixelout<=1'b1;
4224: pixelout<=1'b1;
4225: pixelout<=1'b1;
4226: pixelout<=1'b1;
4227: pixelout<=1'b1;
4228: pixelout<=1'b1;
4229: pixelout<=1'b1;
4230: pixelout<=1'b1;
4231: pixelout<=1'b0;
4232: pixelout<=1'b1;
4233: pixelout<=1'b0;
4234: pixelout<=1'b1;
4235: pixelout<=1'b1;
4236: pixelout<=1'b0;
4237: pixelout<=1'b1;
4238: pixelout<=1'b1;
4239: pixelout<=1'b1;
4240: pixelout<=1'b0;
4241: pixelout<=1'b0;
4242: pixelout<=1'b0;
4243: pixelout<=1'b0;
4244: pixelout<=1'b0;
4245: pixelout<=1'b1;
4246: pixelout<=1'b1;
4247: pixelout<=1'b1;
4248: pixelout<=1'b1;
4249: pixelout<=1'b0;
4250: pixelout<=1'b1;
4251: pixelout<=1'b1;
4252: pixelout<=1'b1;
4253: pixelout<=1'b1;
4254: pixelout<=1'b1;
4255: pixelout<=1'b0;
4256: pixelout<=1'b1;
4257: pixelout<=1'b0;
4258: pixelout<=1'b1;
4259: pixelout<=1'b1;
4260: pixelout<=1'b0;
4261: pixelout<=1'b1;
4262: pixelout<=1'b1;
4263: pixelout<=1'b1;
4264: pixelout<=1'b0;
4265: pixelout<=1'b1;
4266: pixelout<=1'b1;
4267: pixelout<=1'b1;
4268: pixelout<=1'b1;
4269: pixelout<=1'b1;
4270: pixelout<=1'b0;
4271: pixelout<=1'b1;
4272: pixelout<=1'b1;
4273: pixelout<=1'b1;
4274: pixelout<=1'b1;
4275: pixelout<=1'b1;
4276: pixelout<=1'b1;
4277: pixelout<=1'b1;
4278: pixelout<=1'b1;
4279: pixelout<=1'b1;
4280: pixelout<=1'b1;
4281: pixelout<=1'b1;
4282: pixelout<=1'b1;
4283: pixelout<=1'b1;
4284: pixelout<=1'b1;
4285: pixelout<=1'b1;
4286: pixelout<=1'b1;
4287: pixelout<=1'b1;
4288: pixelout<=1'b1;
4289: pixelout<=1'b0;
4290: pixelout<=1'b1;
4291: pixelout<=1'b0;
4292: pixelout<=1'b1;
4293: pixelout<=1'b1;
4294: pixelout<=1'b1;
4295: pixelout<=1'b1;
4296: pixelout<=1'b1;
4297: pixelout<=1'b1;
4298: pixelout<=1'b1;
4299: pixelout<=1'b1;
4300: pixelout<=1'b1;
4301: pixelout<=1'b1;
4302: pixelout<=1'b0;
4303: pixelout<=1'b1;
4304: pixelout<=1'b1;
4305: pixelout<=1'b1;
4306: pixelout<=1'b1;
4307: pixelout<=1'b1;
4308: pixelout<=1'b1;
4309: pixelout<=1'b1;
4310: pixelout<=1'b1;
4311: pixelout<=1'b1;
4312: pixelout<=1'b1;
4313: pixelout<=1'b1;
4314: pixelout<=1'b1;
4315: pixelout<=1'b1;
4316: pixelout<=1'b1;
4317: pixelout<=1'b1;
4318: pixelout<=1'b1;
4319: pixelout<=1'b1;
4320: pixelout<=1'b1;
4321: pixelout<=1'b1;
4322: pixelout<=1'b1;
4323: pixelout<=1'b1;
4324: pixelout<=1'b1;
4325: pixelout<=1'b1;
4326: pixelout<=1'b1;
4327: pixelout<=1'b1;
4328: pixelout<=1'b1;
4329: pixelout<=1'b1;
4330: pixelout<=1'b1;
4331: pixelout<=1'b1;
4332: pixelout<=1'b1;
4333: pixelout<=1'b1;
4334: pixelout<=1'b1;
4335: pixelout<=1'b0;
4336: pixelout<=1'b1;
4337: pixelout<=1'b1;
4338: pixelout<=1'b1;
4339: pixelout<=1'b1;
4340: pixelout<=1'b1;
4341: pixelout<=1'b1;
4342: pixelout<=1'b1;
4343: pixelout<=1'b1;
4344: pixelout<=1'b0;
4345: pixelout<=1'b1;
4346: pixelout<=1'b1;
4347: pixelout<=1'b0;
4348: pixelout<=1'b1;
4349: pixelout<=1'b1;
4350: pixelout<=1'b1;
4351: pixelout<=1'b0;
4352: pixelout<=1'b1;
4353: pixelout<=1'b1;
4354: pixelout<=1'b0;
4355: pixelout<=1'b1;
4356: pixelout<=1'b1;
4357: pixelout<=1'b1;
4358: pixelout<=1'b0;
4359: pixelout<=1'b1;
4360: pixelout<=1'b1;
4361: pixelout<=1'b0;
4362: pixelout<=1'b1;
4363: pixelout<=1'b1;
4364: pixelout<=1'b1;
4365: pixelout<=1'b0;
4366: pixelout<=1'b1;
4367: pixelout<=1'b1;
4368: pixelout<=1'b1;
4369: pixelout<=1'b1;
4370: pixelout<=1'b1;
4371: pixelout<=1'b1;
4372: pixelout<=1'b1;
4373: pixelout<=1'b1;
4374: pixelout<=1'b1;
4375: pixelout<=1'b1;
4376: pixelout<=1'b0;
4377: pixelout<=1'b1;
4378: pixelout<=1'b1;
4379: pixelout<=1'b1;
4380: pixelout<=1'b1;
4381: pixelout<=1'b1;
4382: pixelout<=1'b0;
4383: pixelout<=1'b1;
4384: pixelout<=1'b1;
4385: pixelout<=1'b1;
4386: pixelout<=1'b1;
4387: pixelout<=1'b1;
4388: pixelout<=1'b1;
4389: pixelout<=1'b1;
4390: pixelout<=1'b1;
4391: pixelout<=1'b1;
4392: pixelout<=1'b0;
4393: pixelout<=1'b1;
4394: pixelout<=1'b0;
4395: pixelout<=1'b1;
4396: pixelout<=1'b1;
4397: pixelout<=1'b1;
4398: pixelout<=1'b0;
4399: pixelout<=1'b1;
4400: pixelout<=1'b0;
4401: pixelout<=1'b1;
4402: pixelout<=1'b1;
4403: pixelout<=1'b1;
4404: pixelout<=1'b1;
4405: pixelout<=1'b0;
4406: pixelout<=1'b1;
4407: pixelout<=1'b1;
4408: pixelout<=1'b1;
4409: pixelout<=1'b1;
4410: pixelout<=1'b1;
4411: pixelout<=1'b1;
4412: pixelout<=1'b1;
4413: pixelout<=1'b1;
4414: pixelout<=1'b1;
4415: pixelout<=1'b1;
4416: pixelout<=1'b1;
4417: pixelout<=1'b1;
4418: pixelout<=1'b0;
4419: pixelout<=1'b0;
4420: pixelout<=1'b1;
4421: pixelout<=1'b1;
4422: pixelout<=1'b1;
4423: pixelout<=1'b1;
4424: pixelout<=1'b1;
4425: pixelout<=1'b1;
4426: pixelout<=1'b1;
4427: pixelout<=1'b1;
4428: pixelout<=1'b0;
4429: pixelout<=1'b1;
4430: pixelout<=1'b1;
4431: pixelout<=1'b1;
4432: pixelout<=1'b0;
4433: pixelout<=1'b1;
4434: pixelout<=1'b1;
4435: pixelout<=1'b1;
4436: pixelout<=1'b1;
4437: pixelout<=1'b1;
4438: pixelout<=1'b1;
4439: pixelout<=1'b1;
4440: pixelout<=1'b1;
4441: pixelout<=1'b1;
4442: pixelout<=1'b0;
4443: pixelout<=1'b1;
4444: pixelout<=1'b1;
4445: pixelout<=1'b1;
4446: pixelout<=1'b1;
4447: pixelout<=1'b0;
4448: pixelout<=1'b1;
4449: pixelout<=1'b1;
4450: pixelout<=1'b1;
4451: pixelout<=1'b0;
4452: pixelout<=1'b1;
4453: pixelout<=1'b0;
4454: pixelout<=1'b0;
4455: pixelout<=1'b0;
4456: pixelout<=1'b0;
4457: pixelout<=1'b0;
4458: pixelout<=1'b1;
4459: pixelout<=1'b1;
4460: pixelout<=1'b0;
4461: pixelout<=1'b1;
4462: pixelout<=1'b1;
4463: pixelout<=1'b1;
4464: pixelout<=1'b1;
4465: pixelout<=1'b1;
4466: pixelout<=1'b1;
4467: pixelout<=1'b1;
4468: pixelout<=1'b1;
4469: pixelout<=1'b1;
4470: pixelout<=1'b1;
4471: pixelout<=1'b0;
4472: pixelout<=1'b1;
4473: pixelout<=1'b0;
4474: pixelout<=1'b1;
4475: pixelout<=1'b1;
4476: pixelout<=1'b0;
4477: pixelout<=1'b1;
4478: pixelout<=1'b1;
4479: pixelout<=1'b1;
4480: pixelout<=1'b0;
4481: pixelout<=1'b1;
4482: pixelout<=1'b1;
4483: pixelout<=1'b1;
4484: pixelout<=1'b1;
4485: pixelout<=1'b1;
4486: pixelout<=1'b1;
4487: pixelout<=1'b1;
4488: pixelout<=1'b1;
4489: pixelout<=1'b0;
4490: pixelout<=1'b1;
4491: pixelout<=1'b1;
4492: pixelout<=1'b1;
4493: pixelout<=1'b1;
4494: pixelout<=1'b1;
4495: pixelout<=1'b0;
4496: pixelout<=1'b1;
4497: pixelout<=1'b0;
4498: pixelout<=1'b1;
4499: pixelout<=1'b1;
4500: pixelout<=1'b0;
4501: pixelout<=1'b1;
4502: pixelout<=1'b1;
4503: pixelout<=1'b1;
4504: pixelout<=1'b0;
4505: pixelout<=1'b1;
4506: pixelout<=1'b1;
4507: pixelout<=1'b1;
4508: pixelout<=1'b1;
4509: pixelout<=1'b1;
4510: pixelout<=1'b0;
4511: pixelout<=1'b1;
4512: pixelout<=1'b1;
4513: pixelout<=1'b1;
4514: pixelout<=1'b1;
4515: pixelout<=1'b1;
4516: pixelout<=1'b1;
4517: pixelout<=1'b1;
4518: pixelout<=1'b1;
4519: pixelout<=1'b1;
4520: pixelout<=1'b1;
4521: pixelout<=1'b1;
4522: pixelout<=1'b1;
4523: pixelout<=1'b1;
4524: pixelout<=1'b1;
4525: pixelout<=1'b1;
4526: pixelout<=1'b1;
4527: pixelout<=1'b1;
4528: pixelout<=1'b1;
4529: pixelout<=1'b0;
4530: pixelout<=1'b1;
4531: pixelout<=1'b0;
4532: pixelout<=1'b1;
4533: pixelout<=1'b1;
4534: pixelout<=1'b1;
4535: pixelout<=1'b1;
4536: pixelout<=1'b1;
4537: pixelout<=1'b1;
4538: pixelout<=1'b1;
4539: pixelout<=1'b1;
4540: pixelout<=1'b1;
4541: pixelout<=1'b1;
4542: pixelout<=1'b0;
4543: pixelout<=1'b1;
4544: pixelout<=1'b1;
4545: pixelout<=1'b1;
4546: pixelout<=1'b1;
4547: pixelout<=1'b1;
4548: pixelout<=1'b1;
4549: pixelout<=1'b1;
4550: pixelout<=1'b1;
4551: pixelout<=1'b1;
4552: pixelout<=1'b1;
4553: pixelout<=1'b1;
4554: pixelout<=1'b1;
4555: pixelout<=1'b1;
4556: pixelout<=1'b1;
4557: pixelout<=1'b1;
4558: pixelout<=1'b1;
4559: pixelout<=1'b1;
4560: pixelout<=1'b1;
4561: pixelout<=1'b1;
4562: pixelout<=1'b1;
4563: pixelout<=1'b1;
4564: pixelout<=1'b1;
4565: pixelout<=1'b1;
4566: pixelout<=1'b1;
4567: pixelout<=1'b1;
4568: pixelout<=1'b1;
4569: pixelout<=1'b1;
4570: pixelout<=1'b1;
4571: pixelout<=1'b1;
4572: pixelout<=1'b1;
4573: pixelout<=1'b1;
4574: pixelout<=1'b0;
4575: pixelout<=1'b1;
4576: pixelout<=1'b1;
4577: pixelout<=1'b1;
4578: pixelout<=1'b1;
4579: pixelout<=1'b1;
4580: pixelout<=1'b1;
4581: pixelout<=1'b1;
4582: pixelout<=1'b1;
4583: pixelout<=1'b1;
4584: pixelout<=1'b0;
4585: pixelout<=1'b1;
4586: pixelout<=1'b1;
4587: pixelout<=1'b0;
4588: pixelout<=1'b1;
4589: pixelout<=1'b1;
4590: pixelout<=1'b1;
4591: pixelout<=1'b0;
4592: pixelout<=1'b1;
4593: pixelout<=1'b1;
4594: pixelout<=1'b0;
4595: pixelout<=1'b1;
4596: pixelout<=1'b1;
4597: pixelout<=1'b1;
4598: pixelout<=1'b0;
4599: pixelout<=1'b1;
4600: pixelout<=1'b1;
4601: pixelout<=1'b0;
4602: pixelout<=1'b1;
4603: pixelout<=1'b1;
4604: pixelout<=1'b1;
4605: pixelout<=1'b0;
4606: pixelout<=1'b1;
4607: pixelout<=1'b1;
4608: pixelout<=1'b1;
4609: pixelout<=1'b1;
4610: pixelout<=1'b1;
4611: pixelout<=1'b1;
4612: pixelout<=1'b1;
4613: pixelout<=1'b1;
4614: pixelout<=1'b1;
4615: pixelout<=1'b1;
4616: pixelout<=1'b0;
4617: pixelout<=1'b1;
4618: pixelout<=1'b1;
4619: pixelout<=1'b1;
4620: pixelout<=1'b0;
4621: pixelout<=1'b1;
4622: pixelout<=1'b0;
4623: pixelout<=1'b1;
4624: pixelout<=1'b1;
4625: pixelout<=1'b1;
4626: pixelout<=1'b1;
4627: pixelout<=1'b1;
4628: pixelout<=1'b1;
4629: pixelout<=1'b1;
4630: pixelout<=1'b1;
4631: pixelout<=1'b1;
4632: pixelout<=1'b0;
4633: pixelout<=1'b1;
4634: pixelout<=1'b0;
4635: pixelout<=1'b1;
4636: pixelout<=1'b1;
4637: pixelout<=1'b1;
4638: pixelout<=1'b0;
4639: pixelout<=1'b1;
4640: pixelout<=1'b0;
4641: pixelout<=1'b1;
4642: pixelout<=1'b1;
4643: pixelout<=1'b1;
4644: pixelout<=1'b1;
4645: pixelout<=1'b0;
4646: pixelout<=1'b1;
4647: pixelout<=1'b1;
4648: pixelout<=1'b0;
4649: pixelout<=1'b0;
4650: pixelout<=1'b1;
4651: pixelout<=1'b1;
4652: pixelout<=1'b1;
4653: pixelout<=1'b1;
4654: pixelout<=1'b1;
4655: pixelout<=1'b1;
4656: pixelout<=1'b1;
4657: pixelout<=1'b1;
4658: pixelout<=1'b1;
4659: pixelout<=1'b1;
4660: pixelout<=1'b0;
4661: pixelout<=1'b1;
4662: pixelout<=1'b0;
4663: pixelout<=1'b1;
4664: pixelout<=1'b1;
4665: pixelout<=1'b1;
4666: pixelout<=1'b1;
4667: pixelout<=1'b1;
4668: pixelout<=1'b0;
4669: pixelout<=1'b1;
4670: pixelout<=1'b1;
4671: pixelout<=1'b1;
4672: pixelout<=1'b0;
4673: pixelout<=1'b1;
4674: pixelout<=1'b1;
4675: pixelout<=1'b1;
4676: pixelout<=1'b1;
4677: pixelout<=1'b1;
4678: pixelout<=1'b1;
4679: pixelout<=1'b1;
4680: pixelout<=1'b1;
4681: pixelout<=1'b1;
4682: pixelout<=1'b0;
4683: pixelout<=1'b1;
4684: pixelout<=1'b1;
4685: pixelout<=1'b1;
4686: pixelout<=1'b1;
4687: pixelout<=1'b0;
4688: pixelout<=1'b1;
4689: pixelout<=1'b1;
4690: pixelout<=1'b1;
4691: pixelout<=1'b0;
4692: pixelout<=1'b1;
4693: pixelout<=1'b0;
4694: pixelout<=1'b1;
4695: pixelout<=1'b1;
4696: pixelout<=1'b1;
4697: pixelout<=1'b1;
4698: pixelout<=1'b1;
4699: pixelout<=1'b1;
4700: pixelout<=1'b0;
4701: pixelout<=1'b1;
4702: pixelout<=1'b1;
4703: pixelout<=1'b1;
4704: pixelout<=1'b1;
4705: pixelout<=1'b1;
4706: pixelout<=1'b1;
4707: pixelout<=1'b1;
4708: pixelout<=1'b1;
4709: pixelout<=1'b1;
4710: pixelout<=1'b0;
4711: pixelout<=1'b0;
4712: pixelout<=1'b1;
4713: pixelout<=1'b0;
4714: pixelout<=1'b1;
4715: pixelout<=1'b1;
4716: pixelout<=1'b0;
4717: pixelout<=1'b1;
4718: pixelout<=1'b1;
4719: pixelout<=1'b1;
4720: pixelout<=1'b0;
4721: pixelout<=1'b1;
4722: pixelout<=1'b1;
4723: pixelout<=1'b1;
4724: pixelout<=1'b1;
4725: pixelout<=1'b1;
4726: pixelout<=1'b1;
4727: pixelout<=1'b1;
4728: pixelout<=1'b1;
4729: pixelout<=1'b1;
4730: pixelout<=1'b1;
4731: pixelout<=1'b1;
4732: pixelout<=1'b1;
4733: pixelout<=1'b1;
4734: pixelout<=1'b1;
4735: pixelout<=1'b0;
4736: pixelout<=1'b1;
4737: pixelout<=1'b0;
4738: pixelout<=1'b1;
4739: pixelout<=1'b1;
4740: pixelout<=1'b0;
4741: pixelout<=1'b1;
4742: pixelout<=1'b1;
4743: pixelout<=1'b1;
4744: pixelout<=1'b0;
4745: pixelout<=1'b1;
4746: pixelout<=1'b1;
4747: pixelout<=1'b1;
4748: pixelout<=1'b1;
4749: pixelout<=1'b1;
4750: pixelout<=1'b0;
4751: pixelout<=1'b1;
4752: pixelout<=1'b1;
4753: pixelout<=1'b1;
4754: pixelout<=1'b1;
4755: pixelout<=1'b1;
4756: pixelout<=1'b1;
4757: pixelout<=1'b1;
4758: pixelout<=1'b1;
4759: pixelout<=1'b1;
4760: pixelout<=1'b1;
4761: pixelout<=1'b1;
4762: pixelout<=1'b1;
4763: pixelout<=1'b1;
4764: pixelout<=1'b1;
4765: pixelout<=1'b0;
4766: pixelout<=1'b1;
4767: pixelout<=1'b1;
4768: pixelout<=1'b1;
4769: pixelout<=1'b0;
4770: pixelout<=1'b1;
4771: pixelout<=1'b0;
4772: pixelout<=1'b1;
4773: pixelout<=1'b1;
4774: pixelout<=1'b1;
4775: pixelout<=1'b1;
4776: pixelout<=1'b1;
4777: pixelout<=1'b1;
4778: pixelout<=1'b1;
4779: pixelout<=1'b1;
4780: pixelout<=1'b1;
4781: pixelout<=1'b1;
4782: pixelout<=1'b0;
4783: pixelout<=1'b1;
4784: pixelout<=1'b1;
4785: pixelout<=1'b1;
4786: pixelout<=1'b1;
4787: pixelout<=1'b1;
4788: pixelout<=1'b1;
4789: pixelout<=1'b1;
4790: pixelout<=1'b1;
4791: pixelout<=1'b1;
4792: pixelout<=1'b1;
4793: pixelout<=1'b1;
4794: pixelout<=1'b1;
4795: pixelout<=1'b1;
4796: pixelout<=1'b1;
4797: pixelout<=1'b1;
4798: pixelout<=1'b1;
4799: pixelout<=1'b1;
4800: pixelout<=1'b1;
4801: pixelout<=1'b1;
4802: pixelout<=1'b1;
4803: pixelout<=1'b1;
4804: pixelout<=1'b1;
4805: pixelout<=1'b1;
4806: pixelout<=1'b1;
4807: pixelout<=1'b1;
4808: pixelout<=1'b1;
4809: pixelout<=1'b1;
4810: pixelout<=1'b1;
4811: pixelout<=1'b1;
4812: pixelout<=1'b1;
4813: pixelout<=1'b1;
4814: pixelout<=1'b0;
4815: pixelout<=1'b0;
4816: pixelout<=1'b0;
4817: pixelout<=1'b0;
4818: pixelout<=1'b0;
4819: pixelout<=1'b1;
4820: pixelout<=1'b1;
4821: pixelout<=1'b1;
4822: pixelout<=1'b0;
4823: pixelout<=1'b0;
4824: pixelout<=1'b1;
4825: pixelout<=1'b0;
4826: pixelout<=1'b1;
4827: pixelout<=1'b1;
4828: pixelout<=1'b0;
4829: pixelout<=1'b0;
4830: pixelout<=1'b0;
4831: pixelout<=1'b1;
4832: pixelout<=1'b1;
4833: pixelout<=1'b1;
4834: pixelout<=1'b0;
4835: pixelout<=1'b1;
4836: pixelout<=1'b1;
4837: pixelout<=1'b1;
4838: pixelout<=1'b1;
4839: pixelout<=1'b0;
4840: pixelout<=1'b0;
4841: pixelout<=1'b1;
4842: pixelout<=1'b1;
4843: pixelout<=1'b1;
4844: pixelout<=1'b1;
4845: pixelout<=1'b1;
4846: pixelout<=1'b1;
4847: pixelout<=1'b1;
4848: pixelout<=1'b1;
4849: pixelout<=1'b1;
4850: pixelout<=1'b1;
4851: pixelout<=1'b1;
4852: pixelout<=1'b1;
4853: pixelout<=1'b1;
4854: pixelout<=1'b1;
4855: pixelout<=1'b1;
4856: pixelout<=1'b1;
4857: pixelout<=1'b0;
4858: pixelout<=1'b0;
4859: pixelout<=1'b0;
4860: pixelout<=1'b1;
4861: pixelout<=1'b1;
4862: pixelout<=1'b1;
4863: pixelout<=1'b0;
4864: pixelout<=1'b0;
4865: pixelout<=1'b0;
4866: pixelout<=1'b1;
4867: pixelout<=1'b1;
4868: pixelout<=1'b1;
4869: pixelout<=1'b1;
4870: pixelout<=1'b1;
4871: pixelout<=1'b1;
4872: pixelout<=1'b0;
4873: pixelout<=1'b1;
4874: pixelout<=1'b1;
4875: pixelout<=1'b0;
4876: pixelout<=1'b0;
4877: pixelout<=1'b0;
4878: pixelout<=1'b0;
4879: pixelout<=1'b1;
4880: pixelout<=1'b0;
4881: pixelout<=1'b1;
4882: pixelout<=1'b1;
4883: pixelout<=1'b1;
4884: pixelout<=1'b1;
4885: pixelout<=1'b1;
4886: pixelout<=1'b0;
4887: pixelout<=1'b0;
4888: pixelout<=1'b1;
4889: pixelout<=1'b1;
4890: pixelout<=1'b1;
4891: pixelout<=1'b1;
4892: pixelout<=1'b1;
4893: pixelout<=1'b0;
4894: pixelout<=1'b0;
4895: pixelout<=1'b0;
4896: pixelout<=1'b1;
4897: pixelout<=1'b0;
4898: pixelout<=1'b0;
4899: pixelout<=1'b0;
4900: pixelout<=1'b0;
4901: pixelout<=1'b1;
4902: pixelout<=1'b0;
4903: pixelout<=1'b1;
4904: pixelout<=1'b1;
4905: pixelout<=1'b1;
4906: pixelout<=1'b1;
4907: pixelout<=1'b1;
4908: pixelout<=1'b0;
4909: pixelout<=1'b1;
4910: pixelout<=1'b1;
4911: pixelout<=1'b1;
4912: pixelout<=1'b1;
4913: pixelout<=1'b0;
4914: pixelout<=1'b0;
4915: pixelout<=1'b0;
4916: pixelout<=1'b1;
4917: pixelout<=1'b1;
4918: pixelout<=1'b1;
4919: pixelout<=1'b1;
4920: pixelout<=1'b0;
4921: pixelout<=1'b0;
4922: pixelout<=1'b1;
4923: pixelout<=1'b0;
4924: pixelout<=1'b1;
4925: pixelout<=1'b1;
4926: pixelout<=1'b1;
4927: pixelout<=1'b1;
4928: pixelout<=1'b0;
4929: pixelout<=1'b0;
4930: pixelout<=1'b0;
4931: pixelout<=1'b0;
4932: pixelout<=1'b1;
4933: pixelout<=1'b1;
4934: pixelout<=1'b0;
4935: pixelout<=1'b0;
4936: pixelout<=1'b0;
4937: pixelout<=1'b0;
4938: pixelout<=1'b1;
4939: pixelout<=1'b1;
4940: pixelout<=1'b0;
4941: pixelout<=1'b0;
4942: pixelout<=1'b0;
4943: pixelout<=1'b1;
4944: pixelout<=1'b1;
4945: pixelout<=1'b1;
4946: pixelout<=1'b1;
4947: pixelout<=1'b1;
4948: pixelout<=1'b0;
4949: pixelout<=1'b0;
4950: pixelout<=1'b1;
4951: pixelout<=1'b0;
4952: pixelout<=1'b1;
4953: pixelout<=1'b0;
4954: pixelout<=1'b1;
4955: pixelout<=1'b1;
4956: pixelout<=1'b0;
4957: pixelout<=1'b1;
4958: pixelout<=1'b1;
4959: pixelout<=1'b1;
4960: pixelout<=1'b0;
4961: pixelout<=1'b1;
4962: pixelout<=1'b1;
4963: pixelout<=1'b1;
4964: pixelout<=1'b1;
4965: pixelout<=1'b1;
4966: pixelout<=1'b1;
4967: pixelout<=1'b1;
4968: pixelout<=1'b1;
4969: pixelout<=1'b1;
4970: pixelout<=1'b1;
4971: pixelout<=1'b1;
4972: pixelout<=1'b1;
4973: pixelout<=1'b1;
4974: pixelout<=1'b1;
4975: pixelout<=1'b0;
4976: pixelout<=1'b1;
4977: pixelout<=1'b0;
4978: pixelout<=1'b1;
4979: pixelout<=1'b1;
4980: pixelout<=1'b0;
4981: pixelout<=1'b1;
4982: pixelout<=1'b1;
4983: pixelout<=1'b1;
4984: pixelout<=1'b0;
4985: pixelout<=1'b0;
4986: pixelout<=1'b0;
4987: pixelout<=1'b0;
4988: pixelout<=1'b0;
4989: pixelout<=1'b1;
4990: pixelout<=1'b1;
4991: pixelout<=1'b0;
4992: pixelout<=1'b0;
4993: pixelout<=1'b0;
4994: pixelout<=1'b1;
4995: pixelout<=1'b1;
4996: pixelout<=1'b1;
4997: pixelout<=1'b0;
4998: pixelout<=1'b0;
4999: pixelout<=1'b0;
5000: pixelout<=1'b0;
5001: pixelout<=1'b0;
5002: pixelout<=1'b1;
5003: pixelout<=1'b1;
5004: pixelout<=1'b1;
5005: pixelout<=1'b1;
5006: pixelout<=1'b0;
5007: pixelout<=1'b0;
5008: pixelout<=1'b0;
5009: pixelout<=1'b1;
5010: pixelout<=1'b1;
5011: pixelout<=1'b1;
5012: pixelout<=1'b0;
5013: pixelout<=1'b0;
5014: pixelout<=1'b0;
5015: pixelout<=1'b1;
5016: pixelout<=1'b1;
5017: pixelout<=1'b1;
5018: pixelout<=1'b1;
5019: pixelout<=1'b0;
5020: pixelout<=1'b0;
5021: pixelout<=1'b0;
5022: pixelout<=1'b1;
5023: pixelout<=1'b1;
5024: pixelout<=1'b1;
5025: pixelout<=1'b1;
5026: pixelout<=1'b1;
5027: pixelout<=1'b1;
5028: pixelout<=1'b1;
5029: pixelout<=1'b1;
5030: pixelout<=1'b1;
5031: pixelout<=1'b1;
5032: pixelout<=1'b1;
5033: pixelout<=1'b1;
5034: pixelout<=1'b1;
5035: pixelout<=1'b1;
5036: pixelout<=1'b1;
5037: pixelout<=1'b1;
5038: pixelout<=1'b1;
5039: pixelout<=1'b1;
5040: pixelout<=1'b1;
5041: pixelout<=1'b1;
5042: pixelout<=1'b1;
5043: pixelout<=1'b1;
5044: pixelout<=1'b1;
5045: pixelout<=1'b1;
5046: pixelout<=1'b1;
5047: pixelout<=1'b1;
5048: pixelout<=1'b1;
5049: pixelout<=1'b1;
5050: pixelout<=1'b1;
5051: pixelout<=1'b1;
5052: pixelout<=1'b1;
5053: pixelout<=1'b1;
5054: pixelout<=1'b1;
5055: pixelout<=1'b1;
5056: pixelout<=1'b1;
5057: pixelout<=1'b1;
5058: pixelout<=1'b1;
5059: pixelout<=1'b1;
5060: pixelout<=1'b1;
5061: pixelout<=1'b1;
5062: pixelout<=1'b1;
5063: pixelout<=1'b1;
5064: pixelout<=1'b1;
5065: pixelout<=1'b1;
5066: pixelout<=1'b1;
5067: pixelout<=1'b1;
5068: pixelout<=1'b1;
5069: pixelout<=1'b1;
5070: pixelout<=1'b1;
5071: pixelout<=1'b1;
5072: pixelout<=1'b1;
5073: pixelout<=1'b1;
5074: pixelout<=1'b1;
5075: pixelout<=1'b1;
5076: pixelout<=1'b1;
5077: pixelout<=1'b1;
5078: pixelout<=1'b1;
5079: pixelout<=1'b1;
5080: pixelout<=1'b1;
5081: pixelout<=1'b1;
5082: pixelout<=1'b1;
5083: pixelout<=1'b1;
5084: pixelout<=1'b1;
5085: pixelout<=1'b1;
5086: pixelout<=1'b1;
5087: pixelout<=1'b1;
5088: pixelout<=1'b1;
5089: pixelout<=1'b1;
5090: pixelout<=1'b1;
5091: pixelout<=1'b1;
5092: pixelout<=1'b1;
5093: pixelout<=1'b1;
5094: pixelout<=1'b1;
5095: pixelout<=1'b1;
5096: pixelout<=1'b1;
5097: pixelout<=1'b1;
5098: pixelout<=1'b1;
5099: pixelout<=1'b1;
5100: pixelout<=1'b1;
5101: pixelout<=1'b1;
5102: pixelout<=1'b1;
5103: pixelout<=1'b1;
5104: pixelout<=1'b1;
5105: pixelout<=1'b1;
5106: pixelout<=1'b1;
5107: pixelout<=1'b1;
5108: pixelout<=1'b1;
5109: pixelout<=1'b1;
5110: pixelout<=1'b1;
5111: pixelout<=1'b1;
5112: pixelout<=1'b1;
5113: pixelout<=1'b1;
5114: pixelout<=1'b1;
5115: pixelout<=1'b1;
5116: pixelout<=1'b1;
5117: pixelout<=1'b1;
5118: pixelout<=1'b0;
5119: pixelout<=1'b1;
5120: pixelout<=1'b1;
5121: pixelout<=1'b1;
5122: pixelout<=1'b1;
5123: pixelout<=1'b1;
5124: pixelout<=1'b1;
5125: pixelout<=1'b1;
5126: pixelout<=1'b1;
5127: pixelout<=1'b1;
5128: pixelout<=1'b1;
5129: pixelout<=1'b1;
5130: pixelout<=1'b1;
5131: pixelout<=1'b1;
5132: pixelout<=1'b1;
5133: pixelout<=1'b1;
5134: pixelout<=1'b1;
5135: pixelout<=1'b1;
5136: pixelout<=1'b1;
5137: pixelout<=1'b1;
5138: pixelout<=1'b1;
5139: pixelout<=1'b1;
5140: pixelout<=1'b1;
5141: pixelout<=1'b1;
5142: pixelout<=1'b1;
5143: pixelout<=1'b1;
5144: pixelout<=1'b1;
5145: pixelout<=1'b1;
5146: pixelout<=1'b1;
5147: pixelout<=1'b1;
5148: pixelout<=1'b1;
5149: pixelout<=1'b1;
5150: pixelout<=1'b1;
5151: pixelout<=1'b1;
5152: pixelout<=1'b1;
5153: pixelout<=1'b1;
5154: pixelout<=1'b1;
5155: pixelout<=1'b1;
5156: pixelout<=1'b1;
5157: pixelout<=1'b1;
5158: pixelout<=1'b1;
5159: pixelout<=1'b1;
5160: pixelout<=1'b1;
5161: pixelout<=1'b1;
5162: pixelout<=1'b1;
5163: pixelout<=1'b1;
5164: pixelout<=1'b1;
5165: pixelout<=1'b1;
5166: pixelout<=1'b1;
5167: pixelout<=1'b1;
5168: pixelout<=1'b1;
5169: pixelout<=1'b1;
5170: pixelout<=1'b1;
5171: pixelout<=1'b0;
5172: pixelout<=1'b1;
5173: pixelout<=1'b1;
5174: pixelout<=1'b1;
5175: pixelout<=1'b1;
5176: pixelout<=1'b1;
5177: pixelout<=1'b1;
5178: pixelout<=1'b1;
5179: pixelout<=1'b1;
5180: pixelout<=1'b1;
5181: pixelout<=1'b1;
5182: pixelout<=1'b1;
5183: pixelout<=1'b1;
5184: pixelout<=1'b1;
5185: pixelout<=1'b1;
5186: pixelout<=1'b1;
5187: pixelout<=1'b1;
5188: pixelout<=1'b1;
5189: pixelout<=1'b1;
5190: pixelout<=1'b1;
5191: pixelout<=1'b1;
5192: pixelout<=1'b1;
5193: pixelout<=1'b1;
5194: pixelout<=1'b1;
5195: pixelout<=1'b1;
5196: pixelout<=1'b1;
5197: pixelout<=1'b1;
5198: pixelout<=1'b1;
5199: pixelout<=1'b1;
5200: pixelout<=1'b1;
5201: pixelout<=1'b1;
5202: pixelout<=1'b1;
5203: pixelout<=1'b1;
5204: pixelout<=1'b1;
5205: pixelout<=1'b1;
5206: pixelout<=1'b1;
5207: pixelout<=1'b1;
5208: pixelout<=1'b1;
5209: pixelout<=1'b1;
5210: pixelout<=1'b1;
5211: pixelout<=1'b1;
5212: pixelout<=1'b1;
5213: pixelout<=1'b1;
5214: pixelout<=1'b1;
5215: pixelout<=1'b1;
5216: pixelout<=1'b1;
5217: pixelout<=1'b1;
5218: pixelout<=1'b1;
5219: pixelout<=1'b1;
5220: pixelout<=1'b1;
5221: pixelout<=1'b1;
5222: pixelout<=1'b1;
5223: pixelout<=1'b1;
5224: pixelout<=1'b1;
5225: pixelout<=1'b1;
5226: pixelout<=1'b1;
5227: pixelout<=1'b1;
5228: pixelout<=1'b1;
5229: pixelout<=1'b1;
5230: pixelout<=1'b1;
5231: pixelout<=1'b1;
5232: pixelout<=1'b1;
5233: pixelout<=1'b1;
5234: pixelout<=1'b1;
5235: pixelout<=1'b1;
5236: pixelout<=1'b1;
5237: pixelout<=1'b1;
5238: pixelout<=1'b1;
5239: pixelout<=1'b1;
5240: pixelout<=1'b1;
5241: pixelout<=1'b1;
5242: pixelout<=1'b1;
5243: pixelout<=1'b1;
5244: pixelout<=1'b1;
5245: pixelout<=1'b1;
5246: pixelout<=1'b1;
5247: pixelout<=1'b1;
5248: pixelout<=1'b1;
5249: pixelout<=1'b1;
5250: pixelout<=1'b1;
5251: pixelout<=1'b1;
5252: pixelout<=1'b1;
5253: pixelout<=1'b1;
5254: pixelout<=1'b1;
5255: pixelout<=1'b1;
5256: pixelout<=1'b1;
5257: pixelout<=1'b1;
5258: pixelout<=1'b1;
5259: pixelout<=1'b1;
5260: pixelout<=1'b1;
5261: pixelout<=1'b1;
5262: pixelout<=1'b1;
5263: pixelout<=1'b1;
5264: pixelout<=1'b1;
5265: pixelout<=1'b1;
5266: pixelout<=1'b1;
5267: pixelout<=1'b1;
5268: pixelout<=1'b1;
5269: pixelout<=1'b1;
5270: pixelout<=1'b1;
5271: pixelout<=1'b1;
5272: pixelout<=1'b1;
5273: pixelout<=1'b1;
5274: pixelout<=1'b1;
5275: pixelout<=1'b1;
5276: pixelout<=1'b1;
5277: pixelout<=1'b1;
5278: pixelout<=1'b1;
5279: pixelout<=1'b1;
5280: pixelout<=1'b1;
5281: pixelout<=1'b1;
5282: pixelout<=1'b1;
5283: pixelout<=1'b1;
5284: pixelout<=1'b1;
5285: pixelout<=1'b1;
5286: pixelout<=1'b1;
5287: pixelout<=1'b1;
5288: pixelout<=1'b1;
5289: pixelout<=1'b1;
5290: pixelout<=1'b1;
5291: pixelout<=1'b1;
5292: pixelout<=1'b1;
5293: pixelout<=1'b1;
5294: pixelout<=1'b1;
5295: pixelout<=1'b1;
5296: pixelout<=1'b1;
5297: pixelout<=1'b1;
5298: pixelout<=1'b1;
5299: pixelout<=1'b1;
5300: pixelout<=1'b1;
5301: pixelout<=1'b1;
5302: pixelout<=1'b1;
5303: pixelout<=1'b1;
5304: pixelout<=1'b1;
5305: pixelout<=1'b1;
5306: pixelout<=1'b1;
5307: pixelout<=1'b1;
5308: pixelout<=1'b1;
5309: pixelout<=1'b1;
5310: pixelout<=1'b1;
5311: pixelout<=1'b1;
5312: pixelout<=1'b1;
5313: pixelout<=1'b1;
5314: pixelout<=1'b1;
5315: pixelout<=1'b1;
5316: pixelout<=1'b1;
5317: pixelout<=1'b1;
5318: pixelout<=1'b1;
5319: pixelout<=1'b1;
5320: pixelout<=1'b1;
5321: pixelout<=1'b1;
5322: pixelout<=1'b1;
5323: pixelout<=1'b1;
5324: pixelout<=1'b1;
5325: pixelout<=1'b1;
5326: pixelout<=1'b1;
5327: pixelout<=1'b1;
5328: pixelout<=1'b1;
5329: pixelout<=1'b1;
5330: pixelout<=1'b1;
5331: pixelout<=1'b1;
5332: pixelout<=1'b1;
5333: pixelout<=1'b1;
5334: pixelout<=1'b1;
5335: pixelout<=1'b1;
5336: pixelout<=1'b1;
5337: pixelout<=1'b1;
5338: pixelout<=1'b1;
5339: pixelout<=1'b1;
5340: pixelout<=1'b1;
5341: pixelout<=1'b1;
5342: pixelout<=1'b1;
5343: pixelout<=1'b1;
5344: pixelout<=1'b1;
5345: pixelout<=1'b1;
5346: pixelout<=1'b1;
5347: pixelout<=1'b1;
5348: pixelout<=1'b1;
5349: pixelout<=1'b1;
5350: pixelout<=1'b1;
5351: pixelout<=1'b1;
5352: pixelout<=1'b1;
5353: pixelout<=1'b1;
5354: pixelout<=1'b1;
5355: pixelout<=1'b0;
5356: pixelout<=1'b0;
5357: pixelout<=1'b0;
5358: pixelout<=1'b1;
5359: pixelout<=1'b1;
5360: pixelout<=1'b1;
5361: pixelout<=1'b1;
5362: pixelout<=1'b1;
5363: pixelout<=1'b1;
5364: pixelout<=1'b1;
5365: pixelout<=1'b1;
5366: pixelout<=1'b1;
5367: pixelout<=1'b1;
5368: pixelout<=1'b1;
5369: pixelout<=1'b1;
5370: pixelout<=1'b1;
5371: pixelout<=1'b1;
5372: pixelout<=1'b1;
5373: pixelout<=1'b1;
5374: pixelout<=1'b1;
5375: pixelout<=1'b1;
5376: pixelout<=1'b1;
5377: pixelout<=1'b1;
5378: pixelout<=1'b1;
5379: pixelout<=1'b1;
5380: pixelout<=1'b1;
5381: pixelout<=1'b1;
5382: pixelout<=1'b1;
5383: pixelout<=1'b1;
5384: pixelout<=1'b1;
5385: pixelout<=1'b1;
5386: pixelout<=1'b1;
5387: pixelout<=1'b1;
5388: pixelout<=1'b1;
5389: pixelout<=1'b1;
5390: pixelout<=1'b1;
5391: pixelout<=1'b1;
5392: pixelout<=1'b1;
5393: pixelout<=1'b1;
5394: pixelout<=1'b1;
5395: pixelout<=1'b1;
5396: pixelout<=1'b1;
5397: pixelout<=1'b1;
5398: pixelout<=1'b1;
5399: pixelout<=1'b1;
5400: pixelout<=1'b1;
5401: pixelout<=1'b1;
5402: pixelout<=1'b1;
5403: pixelout<=1'b1;
5404: pixelout<=1'b1;
5405: pixelout<=1'b1;
5406: pixelout<=1'b1;
5407: pixelout<=1'b1;
5408: pixelout<=1'b0;
5409: pixelout<=1'b0;
5410: pixelout<=1'b0;
5411: pixelout<=1'b1;
5412: pixelout<=1'b1;
5413: pixelout<=1'b1;
5414: pixelout<=1'b1;
5415: pixelout<=1'b1;
5416: pixelout<=1'b1;
5417: pixelout<=1'b1;
5418: pixelout<=1'b1;
5419: pixelout<=1'b1;
5420: pixelout<=1'b1;
5421: pixelout<=1'b1;
5422: pixelout<=1'b1;
5423: pixelout<=1'b1;
5424: pixelout<=1'b1;
5425: pixelout<=1'b1;
5426: pixelout<=1'b1;
5427: pixelout<=1'b1;
5428: pixelout<=1'b1;
5429: pixelout<=1'b1;
5430: pixelout<=1'b1;
5431: pixelout<=1'b1;
5432: pixelout<=1'b1;
5433: pixelout<=1'b1;
5434: pixelout<=1'b1;
5435: pixelout<=1'b1;
5436: pixelout<=1'b1;
5437: pixelout<=1'b1;
5438: pixelout<=1'b1;
5439: pixelout<=1'b1;
5440: pixelout<=1'b1;
5441: pixelout<=1'b1;
5442: pixelout<=1'b1;
5443: pixelout<=1'b1;
5444: pixelout<=1'b1;
5445: pixelout<=1'b1;
5446: pixelout<=1'b1;
5447: pixelout<=1'b1;
5448: pixelout<=1'b1;
5449: pixelout<=1'b1;
5450: pixelout<=1'b1;
5451: pixelout<=1'b1;
5452: pixelout<=1'b1;
5453: pixelout<=1'b1;
5454: pixelout<=1'b1;
5455: pixelout<=1'b1;
5456: pixelout<=1'b1;
5457: pixelout<=1'b1;
5458: pixelout<=1'b1;
5459: pixelout<=1'b1;
5460: pixelout<=1'b1;
5461: pixelout<=1'b1;
5462: pixelout<=1'b1;
5463: pixelout<=1'b1;
5464: pixelout<=1'b1;
5465: pixelout<=1'b1;
5466: pixelout<=1'b1;
5467: pixelout<=1'b1;
5468: pixelout<=1'b1;
5469: pixelout<=1'b1;
5470: pixelout<=1'b1;
5471: pixelout<=1'b1;
5472: pixelout<=1'b1;
5473: pixelout<=1'b1;
5474: pixelout<=1'b1;
5475: pixelout<=1'b1;
5476: pixelout<=1'b1;
5477: pixelout<=1'b1;
5478: pixelout<=1'b1;
5479: pixelout<=1'b1;
5480: pixelout<=1'b1;
5481: pixelout<=1'b1;
5482: pixelout<=1'b1;
5483: pixelout<=1'b1;
5484: pixelout<=1'b1;
5485: pixelout<=1'b1;
5486: pixelout<=1'b1;
5487: pixelout<=1'b1;
5488: pixelout<=1'b1;
5489: pixelout<=1'b1;
5490: pixelout<=1'b1;
5491: pixelout<=1'b1;
5492: pixelout<=1'b1;
5493: pixelout<=1'b1;
5494: pixelout<=1'b1;
5495: pixelout<=1'b1;
5496: pixelout<=1'b1;
5497: pixelout<=1'b1;
5498: pixelout<=1'b1;
5499: pixelout<=1'b1;
5500: pixelout<=1'b1;
5501: pixelout<=1'b1;
5502: pixelout<=1'b1;
5503: pixelout<=1'b1;
5504: pixelout<=1'b1;
5505: pixelout<=1'b1;
5506: pixelout<=1'b1;
5507: pixelout<=1'b1;
5508: pixelout<=1'b1;
5509: pixelout<=1'b1;
5510: pixelout<=1'b1;
5511: pixelout<=1'b1;
5512: pixelout<=1'b1;
5513: pixelout<=1'b1;
5514: pixelout<=1'b1;
5515: pixelout<=1'b1;
5516: pixelout<=1'b1;
5517: pixelout<=1'b1;
5518: pixelout<=1'b1;
5519: pixelout<=1'b1;
5520: pixelout<=1'b1;
5521: pixelout<=1'b1;
5522: pixelout<=1'b1;
5523: pixelout<=1'b1;
5524: pixelout<=1'b1;
5525: pixelout<=1'b1;
5526: pixelout<=1'b1;
5527: pixelout<=1'b1;
5528: pixelout<=1'b1;
5529: pixelout<=1'b1;
5530: pixelout<=1'b1;
5531: pixelout<=1'b1;
5532: pixelout<=1'b1;
5533: pixelout<=1'b1;
5534: pixelout<=1'b1;
5535: pixelout<=1'b1;
5536: pixelout<=1'b1;
5537: pixelout<=1'b1;
5538: pixelout<=1'b1;
5539: pixelout<=1'b1;
5540: pixelout<=1'b1;
5541: pixelout<=1'b1;
5542: pixelout<=1'b1;
5543: pixelout<=1'b1;
5544: pixelout<=1'b1;
5545: pixelout<=1'b1;
5546: pixelout<=1'b1;
5547: pixelout<=1'b1;
5548: pixelout<=1'b1;
5549: pixelout<=1'b1;
5550: pixelout<=1'b1;
5551: pixelout<=1'b1;
5552: pixelout<=1'b1;
5553: pixelout<=1'b1;
5554: pixelout<=1'b1;
5555: pixelout<=1'b1;
5556: pixelout<=1'b1;
5557: pixelout<=1'b1;
5558: pixelout<=1'b1;
5559: pixelout<=1'b1;
5560: pixelout<=1'b1;
5561: pixelout<=1'b1;
5562: pixelout<=1'b1;
5563: pixelout<=1'b1;
5564: pixelout<=1'b1;
5565: pixelout<=1'b1;
5566: pixelout<=1'b1;
5567: pixelout<=1'b1;
5568: pixelout<=1'b1;
5569: pixelout<=1'b1;
5570: pixelout<=1'b1;
5571: pixelout<=1'b1;
5572: pixelout<=1'b1;
5573: pixelout<=1'b1;
5574: pixelout<=1'b1;
5575: pixelout<=1'b1;
5576: pixelout<=1'b1;
5577: pixelout<=1'b1;
5578: pixelout<=1'b1;
5579: pixelout<=1'b1;
5580: pixelout<=1'b1;
5581: pixelout<=1'b1;
5582: pixelout<=1'b1;
5583: pixelout<=1'b1;
5584: pixelout<=1'b1;
5585: pixelout<=1'b1;
5586: pixelout<=1'b1;
5587: pixelout<=1'b1;
5588: pixelout<=1'b1;
5589: pixelout<=1'b1;
5590: pixelout<=1'b1;
5591: pixelout<=1'b1;
5592: pixelout<=1'b1;
5593: pixelout<=1'b1;
5594: pixelout<=1'b1;
5595: pixelout<=1'b1;
5596: pixelout<=1'b1;
5597: pixelout<=1'b1;
5598: pixelout<=1'b1;
5599: pixelout<=1'b1;
5600: pixelout<=1'b1;
5601: pixelout<=1'b1;
5602: pixelout<=1'b1;
5603: pixelout<=1'b1;
5604: pixelout<=1'b1;
5605: pixelout<=1'b1;
5606: pixelout<=1'b1;
5607: pixelout<=1'b1;
5608: pixelout<=1'b1;
5609: pixelout<=1'b1;
5610: pixelout<=1'b1;
5611: pixelout<=1'b1;
5612: pixelout<=1'b1;
5613: pixelout<=1'b1;
5614: pixelout<=1'b1;
5615: pixelout<=1'b1;
5616: pixelout<=1'b1;
5617: pixelout<=1'b1;
5618: pixelout<=1'b1;
5619: pixelout<=1'b1;
5620: pixelout<=1'b1;
5621: pixelout<=1'b1;
5622: pixelout<=1'b1;
5623: pixelout<=1'b1;
5624: pixelout<=1'b1;
5625: pixelout<=1'b1;
5626: pixelout<=1'b1;
5627: pixelout<=1'b1;
5628: pixelout<=1'b1;
5629: pixelout<=1'b1;
5630: pixelout<=1'b1;
5631: pixelout<=1'b1;
5632: pixelout<=1'b1;
5633: pixelout<=1'b1;
5634: pixelout<=1'b1;
5635: pixelout<=1'b1;
5636: pixelout<=1'b1;
5637: pixelout<=1'b1;
5638: pixelout<=1'b1;
5639: pixelout<=1'b1;
5640: pixelout<=1'b1;
5641: pixelout<=1'b1;
5642: pixelout<=1'b1;
5643: pixelout<=1'b1;
5644: pixelout<=1'b1;
5645: pixelout<=1'b1;
5646: pixelout<=1'b1;
5647: pixelout<=1'b1;
5648: pixelout<=1'b1;
5649: pixelout<=1'b1;
5650: pixelout<=1'b1;
5651: pixelout<=1'b1;
5652: pixelout<=1'b1;
5653: pixelout<=1'b1;
5654: pixelout<=1'b1;
5655: pixelout<=1'b1;
5656: pixelout<=1'b1;
5657: pixelout<=1'b1;
5658: pixelout<=1'b1;
5659: pixelout<=1'b1;
5660: pixelout<=1'b1;
5661: pixelout<=1'b1;
5662: pixelout<=1'b1;
5663: pixelout<=1'b1;
5664: pixelout<=1'b1;
5665: pixelout<=1'b1;
5666: pixelout<=1'b1;
5667: pixelout<=1'b1;
5668: pixelout<=1'b1;
5669: pixelout<=1'b1;
5670: pixelout<=1'b1;
5671: pixelout<=1'b1;
5672: pixelout<=1'b1;
5673: pixelout<=1'b1;
5674: pixelout<=1'b1;
5675: pixelout<=1'b1;
5676: pixelout<=1'b1;
5677: pixelout<=1'b1;
5678: pixelout<=1'b1;
5679: pixelout<=1'b1;
5680: pixelout<=1'b1;
5681: pixelout<=1'b1;
5682: pixelout<=1'b1;
5683: pixelout<=1'b1;
5684: pixelout<=1'b1;
5685: pixelout<=1'b1;
5686: pixelout<=1'b1;
5687: pixelout<=1'b1;
5688: pixelout<=1'b1;
5689: pixelout<=1'b1;
5690: pixelout<=1'b1;
5691: pixelout<=1'b1;
5692: pixelout<=1'b1;
5693: pixelout<=1'b1;
5694: pixelout<=1'b1;
5695: pixelout<=1'b1;
5696: pixelout<=1'b1;
5697: pixelout<=1'b1;
5698: pixelout<=1'b1;
5699: pixelout<=1'b1;
5700: pixelout<=1'b1;
5701: pixelout<=1'b1;
5702: pixelout<=1'b1;
5703: pixelout<=1'b1;
5704: pixelout<=1'b1;
5705: pixelout<=1'b1;
5706: pixelout<=1'b1;
5707: pixelout<=1'b1;
5708: pixelout<=1'b1;
5709: pixelout<=1'b1;
5710: pixelout<=1'b1;
5711: pixelout<=1'b1;
5712: pixelout<=1'b1;
5713: pixelout<=1'b1;
5714: pixelout<=1'b1;
5715: pixelout<=1'b1;
5716: pixelout<=1'b1;
5717: pixelout<=1'b1;
5718: pixelout<=1'b1;
5719: pixelout<=1'b1;
5720: pixelout<=1'b1;
5721: pixelout<=1'b1;
5722: pixelout<=1'b1;
5723: pixelout<=1'b1;
5724: pixelout<=1'b1;
5725: pixelout<=1'b1;
5726: pixelout<=1'b1;
5727: pixelout<=1'b1;
5728: pixelout<=1'b1;
5729: pixelout<=1'b1;
5730: pixelout<=1'b1;
5731: pixelout<=1'b1;
5732: pixelout<=1'b1;
5733: pixelout<=1'b1;
5734: pixelout<=1'b1;
5735: pixelout<=1'b1;
5736: pixelout<=1'b1;
5737: pixelout<=1'b1;
5738: pixelout<=1'b1;
5739: pixelout<=1'b1;
5740: pixelout<=1'b1;
5741: pixelout<=1'b1;
5742: pixelout<=1'b1;
5743: pixelout<=1'b1;
5744: pixelout<=1'b1;
5745: pixelout<=1'b1;
5746: pixelout<=1'b1;
5747: pixelout<=1'b1;
5748: pixelout<=1'b1;
5749: pixelout<=1'b1;
5750: pixelout<=1'b1;
5751: pixelout<=1'b1;
5752: pixelout<=1'b1;
5753: pixelout<=1'b1;
5754: pixelout<=1'b1;
5755: pixelout<=1'b1;
5756: pixelout<=1'b1;
5757: pixelout<=1'b1;
5758: pixelout<=1'b1;
5759: pixelout<=1'b1;
5760: pixelout<=1'b1;
5761: pixelout<=1'b1;
5762: pixelout<=1'b1;
5763: pixelout<=1'b1;
5764: pixelout<=1'b1;
5765: pixelout<=1'b1;
5766: pixelout<=1'b1;
5767: pixelout<=1'b1;
5768: pixelout<=1'b1;
5769: pixelout<=1'b1;
5770: pixelout<=1'b1;
5771: pixelout<=1'b1;
5772: pixelout<=1'b1;
5773: pixelout<=1'b1;
5774: pixelout<=1'b1;
5775: pixelout<=1'b1;
5776: pixelout<=1'b1;
5777: pixelout<=1'b1;
5778: pixelout<=1'b1;
5779: pixelout<=1'b1;
5780: pixelout<=1'b1;
5781: pixelout<=1'b1;
5782: pixelout<=1'b1;
5783: pixelout<=1'b1;
5784: pixelout<=1'b1;
5785: pixelout<=1'b1;
5786: pixelout<=1'b1;
5787: pixelout<=1'b1;
5788: pixelout<=1'b1;
5789: pixelout<=1'b1;
5790: pixelout<=1'b1;
5791: pixelout<=1'b1;
5792: pixelout<=1'b1;
5793: pixelout<=1'b1;
5794: pixelout<=1'b1;
5795: pixelout<=1'b1;
5796: pixelout<=1'b1;
5797: pixelout<=1'b1;
5798: pixelout<=1'b1;
5799: pixelout<=1'b1;
5800: pixelout<=1'b1;
5801: pixelout<=1'b1;
5802: pixelout<=1'b1;
5803: pixelout<=1'b1;
5804: pixelout<=1'b1;
5805: pixelout<=1'b1;
5806: pixelout<=1'b1;
5807: pixelout<=1'b1;
5808: pixelout<=1'b1;
5809: pixelout<=1'b1;
5810: pixelout<=1'b1;
5811: pixelout<=1'b1;
5812: pixelout<=1'b1;
5813: pixelout<=1'b1;
5814: pixelout<=1'b1;
5815: pixelout<=1'b1;
5816: pixelout<=1'b1;
5817: pixelout<=1'b1;
5818: pixelout<=1'b1;
5819: pixelout<=1'b1;
5820: pixelout<=1'b1;
5821: pixelout<=1'b1;
5822: pixelout<=1'b1;
5823: pixelout<=1'b1;
5824: pixelout<=1'b1;
5825: pixelout<=1'b1;
5826: pixelout<=1'b1;
5827: pixelout<=1'b1;
5828: pixelout<=1'b1;
5829: pixelout<=1'b1;
5830: pixelout<=1'b1;
5831: pixelout<=1'b1;
5832: pixelout<=1'b1;
5833: pixelout<=1'b1;
5834: pixelout<=1'b1;
5835: pixelout<=1'b1;
5836: pixelout<=1'b1;
5837: pixelout<=1'b1;
5838: pixelout<=1'b1;
5839: pixelout<=1'b1;
5840: pixelout<=1'b1;
5841: pixelout<=1'b1;
5842: pixelout<=1'b1;
5843: pixelout<=1'b1;
5844: pixelout<=1'b1;
5845: pixelout<=1'b1;
5846: pixelout<=1'b1;
5847: pixelout<=1'b1;
5848: pixelout<=1'b1;
5849: pixelout<=1'b1;
5850: pixelout<=1'b1;
5851: pixelout<=1'b1;
5852: pixelout<=1'b1;
5853: pixelout<=1'b1;
5854: pixelout<=1'b1;
5855: pixelout<=1'b1;
5856: pixelout<=1'b1;
5857: pixelout<=1'b1;
5858: pixelout<=1'b1;
5859: pixelout<=1'b1;
5860: pixelout<=1'b1;
5861: pixelout<=1'b1;
5862: pixelout<=1'b1;
5863: pixelout<=1'b1;
5864: pixelout<=1'b1;
5865: pixelout<=1'b1;
5866: pixelout<=1'b1;
5867: pixelout<=1'b1;
5868: pixelout<=1'b1;
5869: pixelout<=1'b1;
5870: pixelout<=1'b1;
5871: pixelout<=1'b1;
5872: pixelout<=1'b1;
5873: pixelout<=1'b1;
5874: pixelout<=1'b1;
5875: pixelout<=1'b1;
5876: pixelout<=1'b1;
5877: pixelout<=1'b1;
5878: pixelout<=1'b1;
5879: pixelout<=1'b1;
5880: pixelout<=1'b1;
5881: pixelout<=1'b1;
5882: pixelout<=1'b1;
5883: pixelout<=1'b1;
5884: pixelout<=1'b1;
5885: pixelout<=1'b1;
5886: pixelout<=1'b1;
5887: pixelout<=1'b1;
5888: pixelout<=1'b1;
5889: pixelout<=1'b1;
5890: pixelout<=1'b1;
5891: pixelout<=1'b1;
5892: pixelout<=1'b1;
5893: pixelout<=1'b1;
5894: pixelout<=1'b1;
5895: pixelout<=1'b1;
5896: pixelout<=1'b1;
5897: pixelout<=1'b1;
5898: pixelout<=1'b1;
5899: pixelout<=1'b1;
5900: pixelout<=1'b1;
5901: pixelout<=1'b1;
5902: pixelout<=1'b1;
5903: pixelout<=1'b1;
5904: pixelout<=1'b1;
5905: pixelout<=1'b1;
5906: pixelout<=1'b1;
5907: pixelout<=1'b1;
5908: pixelout<=1'b1;
5909: pixelout<=1'b1;
5910: pixelout<=1'b1;
5911: pixelout<=1'b1;
5912: pixelout<=1'b1;
5913: pixelout<=1'b1;
5914: pixelout<=1'b1;
5915: pixelout<=1'b1;
5916: pixelout<=1'b1;
5917: pixelout<=1'b1;
5918: pixelout<=1'b1;
5919: pixelout<=1'b1;
5920: pixelout<=1'b1;
5921: pixelout<=1'b1;
5922: pixelout<=1'b1;
5923: pixelout<=1'b1;
5924: pixelout<=1'b1;
5925: pixelout<=1'b1;
5926: pixelout<=1'b1;
5927: pixelout<=1'b1;
5928: pixelout<=1'b1;
5929: pixelout<=1'b1;
5930: pixelout<=1'b1;
5931: pixelout<=1'b1;
5932: pixelout<=1'b1;
5933: pixelout<=1'b1;
5934: pixelout<=1'b1;
5935: pixelout<=1'b1;
5936: pixelout<=1'b1;
5937: pixelout<=1'b1;
5938: pixelout<=1'b1;
5939: pixelout<=1'b1;
5940: pixelout<=1'b1;
5941: pixelout<=1'b1;
5942: pixelout<=1'b1;
5943: pixelout<=1'b1;
5944: pixelout<=1'b1;
5945: pixelout<=1'b1;
5946: pixelout<=1'b1;
5947: pixelout<=1'b1;
5948: pixelout<=1'b1;
5949: pixelout<=1'b1;
5950: pixelout<=1'b1;
5951: pixelout<=1'b1;
5952: pixelout<=1'b1;
5953: pixelout<=1'b1;
5954: pixelout<=1'b1;
5955: pixelout<=1'b1;
5956: pixelout<=1'b1;
5957: pixelout<=1'b1;
5958: pixelout<=1'b1;
5959: pixelout<=1'b1;
5960: pixelout<=1'b1;
5961: pixelout<=1'b1;
5962: pixelout<=1'b1;
5963: pixelout<=1'b1;
5964: pixelout<=1'b1;
5965: pixelout<=1'b1;
5966: pixelout<=1'b1;
5967: pixelout<=1'b1;
5968: pixelout<=1'b1;
5969: pixelout<=1'b1;
5970: pixelout<=1'b1;
5971: pixelout<=1'b1;
5972: pixelout<=1'b1;
5973: pixelout<=1'b1;
5974: pixelout<=1'b1;
5975: pixelout<=1'b1;
5976: pixelout<=1'b1;
5977: pixelout<=1'b1;
5978: pixelout<=1'b1;
5979: pixelout<=1'b1;
5980: pixelout<=1'b1;
5981: pixelout<=1'b1;
5982: pixelout<=1'b1;
5983: pixelout<=1'b1;
5984: pixelout<=1'b1;
5985: pixelout<=1'b1;
5986: pixelout<=1'b1;
5987: pixelout<=1'b1;
5988: pixelout<=1'b1;
5989: pixelout<=1'b1;
5990: pixelout<=1'b1;
5991: pixelout<=1'b1;
5992: pixelout<=1'b1;
5993: pixelout<=1'b1;
5994: pixelout<=1'b1;
5995: pixelout<=1'b1;
5996: pixelout<=1'b1;
5997: pixelout<=1'b1;
5998: pixelout<=1'b1;
5999: pixelout<=1'b1;
6000: pixelout<=1'b1;
6001: pixelout<=1'b1;
6002: pixelout<=1'b1;
6003: pixelout<=1'b1;
6004: pixelout<=1'b1;
6005: pixelout<=1'b1;
6006: pixelout<=1'b1;
6007: pixelout<=1'b1;
6008: pixelout<=1'b1;
6009: pixelout<=1'b1;
6010: pixelout<=1'b1;
6011: pixelout<=1'b1;
6012: pixelout<=1'b1;
6013: pixelout<=1'b1;
6014: pixelout<=1'b1;
6015: pixelout<=1'b1;
6016: pixelout<=1'b1;
6017: pixelout<=1'b1;
6018: pixelout<=1'b1;
6019: pixelout<=1'b1;
6020: pixelout<=1'b1;
6021: pixelout<=1'b1;
6022: pixelout<=1'b1;
6023: pixelout<=1'b1;
6024: pixelout<=1'b1;
6025: pixelout<=1'b1;
6026: pixelout<=1'b1;
6027: pixelout<=1'b1;
6028: pixelout<=1'b1;
6029: pixelout<=1'b1;
6030: pixelout<=1'b1;
6031: pixelout<=1'b1;
6032: pixelout<=1'b1;
6033: pixelout<=1'b1;
6034: pixelout<=1'b1;
6035: pixelout<=1'b1;
6036: pixelout<=1'b1;
6037: pixelout<=1'b1;
6038: pixelout<=1'b1;
6039: pixelout<=1'b1;
6040: pixelout<=1'b1;
6041: pixelout<=1'b1;
6042: pixelout<=1'b1;
6043: pixelout<=1'b1;
6044: pixelout<=1'b1;
6045: pixelout<=1'b1;
6046: pixelout<=1'b1;
6047: pixelout<=1'b1;
6048: pixelout<=1'b1;
6049: pixelout<=1'b1;
6050: pixelout<=1'b1;
6051: pixelout<=1'b1;
6052: pixelout<=1'b1;
6053: pixelout<=1'b1;
6054: pixelout<=1'b1;
6055: pixelout<=1'b1;
6056: pixelout<=1'b1;
6057: pixelout<=1'b1;
6058: pixelout<=1'b1;
6059: pixelout<=1'b1;
6060: pixelout<=1'b1;
6061: pixelout<=1'b1;
6062: pixelout<=1'b1;
6063: pixelout<=1'b1;
6064: pixelout<=1'b1;
6065: pixelout<=1'b1;
6066: pixelout<=1'b1;
6067: pixelout<=1'b1;
6068: pixelout<=1'b1;
6069: pixelout<=1'b1;
6070: pixelout<=1'b1;
6071: pixelout<=1'b1;
6072: pixelout<=1'b1;
6073: pixelout<=1'b1;
6074: pixelout<=1'b1;
6075: pixelout<=1'b1;
6076: pixelout<=1'b1;
6077: pixelout<=1'b1;
6078: pixelout<=1'b1;
6079: pixelout<=1'b1;
6080: pixelout<=1'b1;
6081: pixelout<=1'b1;
6082: pixelout<=1'b1;
6083: pixelout<=1'b1;
6084: pixelout<=1'b1;
6085: pixelout<=1'b1;
6086: pixelout<=1'b1;
6087: pixelout<=1'b1;
6088: pixelout<=1'b1;
6089: pixelout<=1'b1;
6090: pixelout<=1'b1;
6091: pixelout<=1'b1;
6092: pixelout<=1'b1;
6093: pixelout<=1'b1;
6094: pixelout<=1'b1;
6095: pixelout<=1'b1;
6096: pixelout<=1'b1;
6097: pixelout<=1'b1;
6098: pixelout<=1'b1;
6099: pixelout<=1'b1;
6100: pixelout<=1'b1;
6101: pixelout<=1'b1;
6102: pixelout<=1'b1;
6103: pixelout<=1'b1;
6104: pixelout<=1'b1;
6105: pixelout<=1'b1;
6106: pixelout<=1'b1;
6107: pixelout<=1'b1;
6108: pixelout<=1'b1;
6109: pixelout<=1'b1;
6110: pixelout<=1'b1;
6111: pixelout<=1'b1;
6112: pixelout<=1'b1;
6113: pixelout<=1'b1;
6114: pixelout<=1'b1;
6115: pixelout<=1'b1;
6116: pixelout<=1'b1;
6117: pixelout<=1'b1;
6118: pixelout<=1'b1;
6119: pixelout<=1'b1;
6120: pixelout<=1'b1;
6121: pixelout<=1'b1;
6122: pixelout<=1'b1;
6123: pixelout<=1'b1;
6124: pixelout<=1'b1;
6125: pixelout<=1'b1;
6126: pixelout<=1'b1;
6127: pixelout<=1'b1;
6128: pixelout<=1'b1;
6129: pixelout<=1'b1;
6130: pixelout<=1'b1;
6131: pixelout<=1'b1;
6132: pixelout<=1'b1;
6133: pixelout<=1'b1;
6134: pixelout<=1'b1;
6135: pixelout<=1'b1;
6136: pixelout<=1'b1;
6137: pixelout<=1'b1;
6138: pixelout<=1'b1;
6139: pixelout<=1'b1;
6140: pixelout<=1'b1;
6141: pixelout<=1'b1;
6142: pixelout<=1'b1;
6143: pixelout<=1'b1;
6144: pixelout<=1'b1;
6145: pixelout<=1'b1;
6146: pixelout<=1'b1;
6147: pixelout<=1'b1;
6148: pixelout<=1'b1;
6149: pixelout<=1'b1;
6150: pixelout<=1'b1;
6151: pixelout<=1'b1;
6152: pixelout<=1'b1;
6153: pixelout<=1'b1;
6154: pixelout<=1'b1;
6155: pixelout<=1'b1;
6156: pixelout<=1'b1;
6157: pixelout<=1'b1;
6158: pixelout<=1'b1;
6159: pixelout<=1'b1;
6160: pixelout<=1'b1;
6161: pixelout<=1'b1;
6162: pixelout<=1'b1;
6163: pixelout<=1'b1;
6164: pixelout<=1'b1;
6165: pixelout<=1'b1;
6166: pixelout<=1'b1;
6167: pixelout<=1'b1;
6168: pixelout<=1'b1;
6169: pixelout<=1'b1;
6170: pixelout<=1'b1;
6171: pixelout<=1'b1;
6172: pixelout<=1'b1;
6173: pixelout<=1'b1;
6174: pixelout<=1'b1;
6175: pixelout<=1'b1;
6176: pixelout<=1'b1;
6177: pixelout<=1'b1;
6178: pixelout<=1'b1;
6179: pixelout<=1'b1;
6180: pixelout<=1'b1;
6181: pixelout<=1'b1;
6182: pixelout<=1'b1;
6183: pixelout<=1'b1;
6184: pixelout<=1'b1;
6185: pixelout<=1'b1;
6186: pixelout<=1'b1;
6187: pixelout<=1'b1;
6188: pixelout<=1'b1;
6189: pixelout<=1'b1;
6190: pixelout<=1'b1;
6191: pixelout<=1'b1;
6192: pixelout<=1'b1;
6193: pixelout<=1'b1;
6194: pixelout<=1'b1;
6195: pixelout<=1'b1;
6196: pixelout<=1'b1;
6197: pixelout<=1'b1;
6198: pixelout<=1'b1;
6199: pixelout<=1'b1;
6200: pixelout<=1'b1;
6201: pixelout<=1'b1;
6202: pixelout<=1'b1;
6203: pixelout<=1'b1;
6204: pixelout<=1'b1;
6205: pixelout<=1'b1;
6206: pixelout<=1'b1;
6207: pixelout<=1'b1;
6208: pixelout<=1'b1;
6209: pixelout<=1'b1;
6210: pixelout<=1'b1;
6211: pixelout<=1'b1;
6212: pixelout<=1'b1;
6213: pixelout<=1'b1;
6214: pixelout<=1'b1;
6215: pixelout<=1'b1;
6216: pixelout<=1'b1;
6217: pixelout<=1'b1;
6218: pixelout<=1'b1;
6219: pixelout<=1'b1;
6220: pixelout<=1'b1;
6221: pixelout<=1'b1;
6222: pixelout<=1'b1;
6223: pixelout<=1'b1;
6224: pixelout<=1'b1;
6225: pixelout<=1'b1;
6226: pixelout<=1'b1;
6227: pixelout<=1'b1;
6228: pixelout<=1'b1;
6229: pixelout<=1'b1;
6230: pixelout<=1'b1;
6231: pixelout<=1'b1;
6232: pixelout<=1'b1;
6233: pixelout<=1'b1;
6234: pixelout<=1'b1;
6235: pixelout<=1'b1;
6236: pixelout<=1'b1;
6237: pixelout<=1'b1;
6238: pixelout<=1'b1;
6239: pixelout<=1'b1;
6240: pixelout<=1'b1;
6241: pixelout<=1'b1;
6242: pixelout<=1'b1;
6243: pixelout<=1'b1;
6244: pixelout<=1'b1;
6245: pixelout<=1'b1;
6246: pixelout<=1'b1;
6247: pixelout<=1'b1;
6248: pixelout<=1'b1;
6249: pixelout<=1'b1;
6250: pixelout<=1'b1;
6251: pixelout<=1'b1;
6252: pixelout<=1'b1;
6253: pixelout<=1'b1;
6254: pixelout<=1'b1;
6255: pixelout<=1'b1;
6256: pixelout<=1'b1;
6257: pixelout<=1'b1;
6258: pixelout<=1'b1;
6259: pixelout<=1'b1;
6260: pixelout<=1'b1;
6261: pixelout<=1'b1;
6262: pixelout<=1'b1;
6263: pixelout<=1'b1;
6264: pixelout<=1'b1;
6265: pixelout<=1'b1;
6266: pixelout<=1'b1;
6267: pixelout<=1'b1;
6268: pixelout<=1'b1;
6269: pixelout<=1'b1;
6270: pixelout<=1'b1;
6271: pixelout<=1'b1;
6272: pixelout<=1'b1;
6273: pixelout<=1'b1;
6274: pixelout<=1'b1;
6275: pixelout<=1'b1;
6276: pixelout<=1'b1;
6277: pixelout<=1'b1;
6278: pixelout<=1'b1;
6279: pixelout<=1'b1;
6280: pixelout<=1'b1;
6281: pixelout<=1'b1;
6282: pixelout<=1'b1;
6283: pixelout<=1'b1;
6284: pixelout<=1'b1;
6285: pixelout<=1'b1;
6286: pixelout<=1'b1;
6287: pixelout<=1'b1;
6288: pixelout<=1'b1;
6289: pixelout<=1'b1;
6290: pixelout<=1'b1;
6291: pixelout<=1'b1;
6292: pixelout<=1'b1;
6293: pixelout<=1'b1;
6294: pixelout<=1'b1;
6295: pixelout<=1'b1;
6296: pixelout<=1'b1;
6297: pixelout<=1'b1;
6298: pixelout<=1'b1;
6299: pixelout<=1'b1;
6300: pixelout<=1'b1;
6301: pixelout<=1'b1;
6302: pixelout<=1'b1;
6303: pixelout<=1'b1;
6304: pixelout<=1'b1;
6305: pixelout<=1'b1;
6306: pixelout<=1'b1;
6307: pixelout<=1'b1;
6308: pixelout<=1'b1;
6309: pixelout<=1'b1;
6310: pixelout<=1'b1;
6311: pixelout<=1'b1;
6312: pixelout<=1'b1;
6313: pixelout<=1'b1;
6314: pixelout<=1'b1;
6315: pixelout<=1'b1;
6316: pixelout<=1'b1;
6317: pixelout<=1'b1;
6318: pixelout<=1'b1;
6319: pixelout<=1'b1;
6320: pixelout<=1'b1;
6321: pixelout<=1'b1;
6322: pixelout<=1'b1;
6323: pixelout<=1'b1;
6324: pixelout<=1'b1;
6325: pixelout<=1'b1;
6326: pixelout<=1'b1;
6327: pixelout<=1'b1;
6328: pixelout<=1'b1;
6329: pixelout<=1'b1;
6330: pixelout<=1'b1;
6331: pixelout<=1'b1;
6332: pixelout<=1'b1;
6333: pixelout<=1'b1;
6334: pixelout<=1'b1;
6335: pixelout<=1'b1;
6336: pixelout<=1'b1;
6337: pixelout<=1'b1;
6338: pixelout<=1'b1;
6339: pixelout<=1'b1;
6340: pixelout<=1'b1;
6341: pixelout<=1'b1;
6342: pixelout<=1'b1;
6343: pixelout<=1'b1;
6344: pixelout<=1'b1;
6345: pixelout<=1'b1;
6346: pixelout<=1'b1;
6347: pixelout<=1'b1;
6348: pixelout<=1'b1;
6349: pixelout<=1'b1;
6350: pixelout<=1'b1;
6351: pixelout<=1'b1;
6352: pixelout<=1'b1;
6353: pixelout<=1'b1;
6354: pixelout<=1'b1;
6355: pixelout<=1'b1;
6356: pixelout<=1'b1;
6357: pixelout<=1'b1;
6358: pixelout<=1'b1;
6359: pixelout<=1'b1;
6360: pixelout<=1'b1;
6361: pixelout<=1'b1;
6362: pixelout<=1'b1;
6363: pixelout<=1'b1;
6364: pixelout<=1'b1;
6365: pixelout<=1'b1;
6366: pixelout<=1'b1;
6367: pixelout<=1'b1;
6368: pixelout<=1'b1;
6369: pixelout<=1'b1;
6370: pixelout<=1'b1;
6371: pixelout<=1'b1;
6372: pixelout<=1'b1;
6373: pixelout<=1'b1;
6374: pixelout<=1'b1;
6375: pixelout<=1'b1;
6376: pixelout<=1'b1;
6377: pixelout<=1'b1;
6378: pixelout<=1'b1;
6379: pixelout<=1'b1;
6380: pixelout<=1'b1;
6381: pixelout<=1'b1;
6382: pixelout<=1'b1;
6383: pixelout<=1'b1;
6384: pixelout<=1'b1;
6385: pixelout<=1'b1;
6386: pixelout<=1'b1;
6387: pixelout<=1'b1;
6388: pixelout<=1'b1;
6389: pixelout<=1'b1;
6390: pixelout<=1'b1;
6391: pixelout<=1'b1;
6392: pixelout<=1'b1;
6393: pixelout<=1'b1;
6394: pixelout<=1'b1;
6395: pixelout<=1'b1;
6396: pixelout<=1'b1;
6397: pixelout<=1'b1;
6398: pixelout<=1'b1;
6399: pixelout<=1'b1;
6400: pixelout<=1'b1;
6401: pixelout<=1'b1;
6402: pixelout<=1'b1;
6403: pixelout<=1'b1;
6404: pixelout<=1'b1;
6405: pixelout<=1'b1;
6406: pixelout<=1'b1;
6407: pixelout<=1'b1;
6408: pixelout<=1'b1;
6409: pixelout<=1'b1;
6410: pixelout<=1'b1;
6411: pixelout<=1'b1;
6412: pixelout<=1'b1;
6413: pixelout<=1'b1;
6414: pixelout<=1'b1;
6415: pixelout<=1'b1;
6416: pixelout<=1'b1;
6417: pixelout<=1'b1;
6418: pixelout<=1'b1;
6419: pixelout<=1'b1;
6420: pixelout<=1'b1;
6421: pixelout<=1'b1;
6422: pixelout<=1'b1;
6423: pixelout<=1'b1;
6424: pixelout<=1'b1;
6425: pixelout<=1'b1;
6426: pixelout<=1'b1;
6427: pixelout<=1'b1;
6428: pixelout<=1'b1;
6429: pixelout<=1'b1;
6430: pixelout<=1'b1;
6431: pixelout<=1'b1;
6432: pixelout<=1'b1;
6433: pixelout<=1'b1;
6434: pixelout<=1'b1;
6435: pixelout<=1'b1;
6436: pixelout<=1'b1;
6437: pixelout<=1'b1;
6438: pixelout<=1'b1;
6439: pixelout<=1'b1;
6440: pixelout<=1'b1;
6441: pixelout<=1'b1;
6442: pixelout<=1'b1;
6443: pixelout<=1'b1;
6444: pixelout<=1'b1;
6445: pixelout<=1'b1;
6446: pixelout<=1'b1;
6447: pixelout<=1'b1;
6448: pixelout<=1'b1;
6449: pixelout<=1'b1;
6450: pixelout<=1'b1;
6451: pixelout<=1'b1;
6452: pixelout<=1'b1;
6453: pixelout<=1'b1;
6454: pixelout<=1'b1;
6455: pixelout<=1'b1;
6456: pixelout<=1'b1;
6457: pixelout<=1'b1;
6458: pixelout<=1'b1;
6459: pixelout<=1'b1;
6460: pixelout<=1'b1;
6461: pixelout<=1'b1;
6462: pixelout<=1'b1;
6463: pixelout<=1'b1;
6464: pixelout<=1'b1;
6465: pixelout<=1'b1;
6466: pixelout<=1'b1;
6467: pixelout<=1'b1;
6468: pixelout<=1'b1;
6469: pixelout<=1'b1;
6470: pixelout<=1'b1;
6471: pixelout<=1'b1;
6472: pixelout<=1'b1;
6473: pixelout<=1'b1;
6474: pixelout<=1'b1;
6475: pixelout<=1'b1;
6476: pixelout<=1'b1;
6477: pixelout<=1'b1;
6478: pixelout<=1'b1;
6479: pixelout<=1'b1;
6480: pixelout<=1'b1;
6481: pixelout<=1'b1;
6482: pixelout<=1'b1;
6483: pixelout<=1'b1;
6484: pixelout<=1'b1;
6485: pixelout<=1'b1;
6486: pixelout<=1'b1;
6487: pixelout<=1'b1;
6488: pixelout<=1'b1;
6489: pixelout<=1'b1;
6490: pixelout<=1'b1;
6491: pixelout<=1'b1;
6492: pixelout<=1'b1;
6493: pixelout<=1'b1;
6494: pixelout<=1'b1;
6495: pixelout<=1'b1;
6496: pixelout<=1'b1;
6497: pixelout<=1'b1;
6498: pixelout<=1'b1;
6499: pixelout<=1'b1;
6500: pixelout<=1'b1;
6501: pixelout<=1'b1;
6502: pixelout<=1'b1;
6503: pixelout<=1'b1;
6504: pixelout<=1'b1;
6505: pixelout<=1'b1;
6506: pixelout<=1'b1;
6507: pixelout<=1'b1;
6508: pixelout<=1'b1;
6509: pixelout<=1'b1;
6510: pixelout<=1'b1;
6511: pixelout<=1'b1;
6512: pixelout<=1'b1;
6513: pixelout<=1'b1;
6514: pixelout<=1'b1;
6515: pixelout<=1'b1;
6516: pixelout<=1'b1;
6517: pixelout<=1'b1;
6518: pixelout<=1'b1;
6519: pixelout<=1'b1;
6520: pixelout<=1'b1;
6521: pixelout<=1'b1;
6522: pixelout<=1'b1;
6523: pixelout<=1'b1;
6524: pixelout<=1'b1;
6525: pixelout<=1'b1;
6526: pixelout<=1'b1;
6527: pixelout<=1'b1;
6528: pixelout<=1'b1;
6529: pixelout<=1'b1;
6530: pixelout<=1'b1;
6531: pixelout<=1'b1;
6532: pixelout<=1'b1;
6533: pixelout<=1'b1;
6534: pixelout<=1'b1;
6535: pixelout<=1'b1;
6536: pixelout<=1'b1;
6537: pixelout<=1'b1;
6538: pixelout<=1'b1;
6539: pixelout<=1'b1;
6540: pixelout<=1'b1;
6541: pixelout<=1'b1;
6542: pixelout<=1'b1;
6543: pixelout<=1'b1;
6544: pixelout<=1'b1;
6545: pixelout<=1'b1;
6546: pixelout<=1'b1;
6547: pixelout<=1'b1;
6548: pixelout<=1'b1;
6549: pixelout<=1'b1;
6550: pixelout<=1'b1;
6551: pixelout<=1'b1;
6552: pixelout<=1'b1;
6553: pixelout<=1'b1;
6554: pixelout<=1'b1;
6555: pixelout<=1'b1;
6556: pixelout<=1'b1;
6557: pixelout<=1'b1;
6558: pixelout<=1'b1;
6559: pixelout<=1'b1;
6560: pixelout<=1'b1;
6561: pixelout<=1'b1;
6562: pixelout<=1'b1;
6563: pixelout<=1'b1;
6564: pixelout<=1'b1;
6565: pixelout<=1'b1;
6566: pixelout<=1'b1;
6567: pixelout<=1'b1;
6568: pixelout<=1'b1;
6569: pixelout<=1'b1;
6570: pixelout<=1'b1;
6571: pixelout<=1'b1;
6572: pixelout<=1'b1;
6573: pixelout<=1'b1;
6574: pixelout<=1'b1;
6575: pixelout<=1'b1;
6576: pixelout<=1'b1;
6577: pixelout<=1'b1;
6578: pixelout<=1'b1;
6579: pixelout<=1'b1;
6580: pixelout<=1'b1;
6581: pixelout<=1'b1;
6582: pixelout<=1'b1;
6583: pixelout<=1'b1;
6584: pixelout<=1'b1;
6585: pixelout<=1'b1;
6586: pixelout<=1'b1;
6587: pixelout<=1'b1;
6588: pixelout<=1'b1;
6589: pixelout<=1'b1;
6590: pixelout<=1'b1;
6591: pixelout<=1'b1;
6592: pixelout<=1'b1;
6593: pixelout<=1'b1;
6594: pixelout<=1'b1;
6595: pixelout<=1'b1;
6596: pixelout<=1'b1;
6597: pixelout<=1'b1;
6598: pixelout<=1'b1;
6599: pixelout<=1'b1;
6600: pixelout<=1'b1;
6601: pixelout<=1'b1;
6602: pixelout<=1'b1;
6603: pixelout<=1'b1;
6604: pixelout<=1'b1;
6605: pixelout<=1'b1;
6606: pixelout<=1'b1;
6607: pixelout<=1'b1;
6608: pixelout<=1'b1;
6609: pixelout<=1'b1;
6610: pixelout<=1'b1;
6611: pixelout<=1'b1;
6612: pixelout<=1'b1;
6613: pixelout<=1'b1;
6614: pixelout<=1'b1;
6615: pixelout<=1'b1;
6616: pixelout<=1'b1;
6617: pixelout<=1'b1;
6618: pixelout<=1'b1;
6619: pixelout<=1'b1;
6620: pixelout<=1'b1;
6621: pixelout<=1'b1;
6622: pixelout<=1'b1;
6623: pixelout<=1'b1;
6624: pixelout<=1'b1;
6625: pixelout<=1'b1;
6626: pixelout<=1'b1;
6627: pixelout<=1'b1;
6628: pixelout<=1'b1;
6629: pixelout<=1'b1;
6630: pixelout<=1'b1;
6631: pixelout<=1'b1;
6632: pixelout<=1'b1;
6633: pixelout<=1'b1;
6634: pixelout<=1'b1;
6635: pixelout<=1'b1;
6636: pixelout<=1'b1;
6637: pixelout<=1'b1;
6638: pixelout<=1'b1;
6639: pixelout<=1'b1;
6640: pixelout<=1'b1;
6641: pixelout<=1'b1;
6642: pixelout<=1'b1;
6643: pixelout<=1'b1;
6644: pixelout<=1'b1;
6645: pixelout<=1'b1;
6646: pixelout<=1'b1;
6647: pixelout<=1'b1;
6648: pixelout<=1'b1;
6649: pixelout<=1'b1;
6650: pixelout<=1'b1;
6651: pixelout<=1'b1;
6652: pixelout<=1'b1;
6653: pixelout<=1'b1;
6654: pixelout<=1'b1;
6655: pixelout<=1'b1;
6656: pixelout<=1'b1;
6657: pixelout<=1'b1;
6658: pixelout<=1'b1;
6659: pixelout<=1'b1;
6660: pixelout<=1'b1;
6661: pixelout<=1'b1;
6662: pixelout<=1'b1;
6663: pixelout<=1'b1;
6664: pixelout<=1'b1;
6665: pixelout<=1'b1;
6666: pixelout<=1'b1;
6667: pixelout<=1'b1;
6668: pixelout<=1'b1;
6669: pixelout<=1'b1;
6670: pixelout<=1'b1;
6671: pixelout<=1'b1;
6672: pixelout<=1'b1;
6673: pixelout<=1'b1;
6674: pixelout<=1'b1;
6675: pixelout<=1'b1;
6676: pixelout<=1'b1;
6677: pixelout<=1'b1;
6678: pixelout<=1'b1;
6679: pixelout<=1'b1;
6680: pixelout<=1'b1;
6681: pixelout<=1'b1;
6682: pixelout<=1'b1;
6683: pixelout<=1'b1;
6684: pixelout<=1'b1;
6685: pixelout<=1'b1;
6686: pixelout<=1'b1;
6687: pixelout<=1'b1;
6688: pixelout<=1'b1;
6689: pixelout<=1'b1;
6690: pixelout<=1'b1;
6691: pixelout<=1'b1;
6692: pixelout<=1'b1;
6693: pixelout<=1'b1;
6694: pixelout<=1'b1;
6695: pixelout<=1'b1;
6696: pixelout<=1'b1;
6697: pixelout<=1'b1;
6698: pixelout<=1'b1;
6699: pixelout<=1'b1;
6700: pixelout<=1'b1;
6701: pixelout<=1'b1;
6702: pixelout<=1'b1;
6703: pixelout<=1'b1;
6704: pixelout<=1'b1;
6705: pixelout<=1'b1;
6706: pixelout<=1'b1;
6707: pixelout<=1'b1;
6708: pixelout<=1'b1;
6709: pixelout<=1'b1;
6710: pixelout<=1'b1;
6711: pixelout<=1'b1;
6712: pixelout<=1'b1;
6713: pixelout<=1'b1;
6714: pixelout<=1'b1;
6715: pixelout<=1'b1;
6716: pixelout<=1'b1;
6717: pixelout<=1'b1;
6718: pixelout<=1'b1;
6719: pixelout<=1'b1;
6720: pixelout<=1'b1;
6721: pixelout<=1'b1;
6722: pixelout<=1'b1;
6723: pixelout<=1'b1;
6724: pixelout<=1'b1;
6725: pixelout<=1'b1;
6726: pixelout<=1'b1;
6727: pixelout<=1'b1;
6728: pixelout<=1'b1;
6729: pixelout<=1'b1;
6730: pixelout<=1'b1;
6731: pixelout<=1'b1;
6732: pixelout<=1'b1;
6733: pixelout<=1'b1;
6734: pixelout<=1'b1;
6735: pixelout<=1'b1;
6736: pixelout<=1'b1;
6737: pixelout<=1'b1;
6738: pixelout<=1'b1;
6739: pixelout<=1'b1;
6740: pixelout<=1'b1;
6741: pixelout<=1'b1;
6742: pixelout<=1'b1;
6743: pixelout<=1'b1;
6744: pixelout<=1'b1;
6745: pixelout<=1'b1;
6746: pixelout<=1'b1;
6747: pixelout<=1'b1;
6748: pixelout<=1'b1;
6749: pixelout<=1'b1;
6750: pixelout<=1'b1;
6751: pixelout<=1'b1;
6752: pixelout<=1'b1;
6753: pixelout<=1'b1;
6754: pixelout<=1'b1;
6755: pixelout<=1'b1;
6756: pixelout<=1'b1;
6757: pixelout<=1'b1;
6758: pixelout<=1'b1;
6759: pixelout<=1'b1;
6760: pixelout<=1'b1;
6761: pixelout<=1'b1;
6762: pixelout<=1'b1;
6763: pixelout<=1'b1;
6764: pixelout<=1'b1;
6765: pixelout<=1'b1;
6766: pixelout<=1'b1;
6767: pixelout<=1'b1;
6768: pixelout<=1'b1;
6769: pixelout<=1'b1;
6770: pixelout<=1'b1;
6771: pixelout<=1'b1;
6772: pixelout<=1'b1;
6773: pixelout<=1'b1;
6774: pixelout<=1'b1;
6775: pixelout<=1'b1;
6776: pixelout<=1'b1;
6777: pixelout<=1'b1;
6778: pixelout<=1'b1;
6779: pixelout<=1'b1;
6780: pixelout<=1'b1;
6781: pixelout<=1'b1;
6782: pixelout<=1'b1;
6783: pixelout<=1'b1;
6784: pixelout<=1'b1;
6785: pixelout<=1'b1;
6786: pixelout<=1'b1;
6787: pixelout<=1'b1;
6788: pixelout<=1'b1;
6789: pixelout<=1'b1;
6790: pixelout<=1'b1;
6791: pixelout<=1'b1;
6792: pixelout<=1'b1;
6793: pixelout<=1'b1;
6794: pixelout<=1'b1;
6795: pixelout<=1'b1;
6796: pixelout<=1'b1;
6797: pixelout<=1'b1;
6798: pixelout<=1'b1;
6799: pixelout<=1'b1;
6800: pixelout<=1'b1;
6801: pixelout<=1'b1;
6802: pixelout<=1'b1;
6803: pixelout<=1'b1;
6804: pixelout<=1'b1;
6805: pixelout<=1'b1;
6806: pixelout<=1'b1;
6807: pixelout<=1'b1;
6808: pixelout<=1'b1;
6809: pixelout<=1'b1;
6810: pixelout<=1'b1;
6811: pixelout<=1'b1;
6812: pixelout<=1'b1;
6813: pixelout<=1'b1;
6814: pixelout<=1'b1;
6815: pixelout<=1'b1;
6816: pixelout<=1'b1;
6817: pixelout<=1'b1;
6818: pixelout<=1'b1;
6819: pixelout<=1'b1;
6820: pixelout<=1'b1;
6821: pixelout<=1'b1;
6822: pixelout<=1'b1;
6823: pixelout<=1'b1;
6824: pixelout<=1'b1;
6825: pixelout<=1'b1;
6826: pixelout<=1'b1;
6827: pixelout<=1'b1;
6828: pixelout<=1'b1;
6829: pixelout<=1'b1;
6830: pixelout<=1'b1;
6831: pixelout<=1'b1;
6832: pixelout<=1'b1;
6833: pixelout<=1'b1;
6834: pixelout<=1'b1;
6835: pixelout<=1'b1;
6836: pixelout<=1'b1;
6837: pixelout<=1'b1;
6838: pixelout<=1'b1;
6839: pixelout<=1'b1;
6840: pixelout<=1'b1;
6841: pixelout<=1'b1;
6842: pixelout<=1'b1;
6843: pixelout<=1'b1;
6844: pixelout<=1'b1;
6845: pixelout<=1'b1;
6846: pixelout<=1'b1;
6847: pixelout<=1'b1;
6848: pixelout<=1'b1;
6849: pixelout<=1'b1;
6850: pixelout<=1'b1;
6851: pixelout<=1'b1;
6852: pixelout<=1'b1;
6853: pixelout<=1'b1;
6854: pixelout<=1'b1;
6855: pixelout<=1'b1;
6856: pixelout<=1'b1;
6857: pixelout<=1'b1;
6858: pixelout<=1'b1;
6859: pixelout<=1'b1;
6860: pixelout<=1'b1;
6861: pixelout<=1'b1;
6862: pixelout<=1'b1;
6863: pixelout<=1'b1;
6864: pixelout<=1'b1;
6865: pixelout<=1'b1;
6866: pixelout<=1'b1;
6867: pixelout<=1'b1;
6868: pixelout<=1'b1;
6869: pixelout<=1'b1;
6870: pixelout<=1'b1;
6871: pixelout<=1'b1;
6872: pixelout<=1'b1;
6873: pixelout<=1'b1;
6874: pixelout<=1'b1;
6875: pixelout<=1'b1;
6876: pixelout<=1'b1;
6877: pixelout<=1'b1;
6878: pixelout<=1'b1;
6879: pixelout<=1'b1;
6880: pixelout<=1'b1;
6881: pixelout<=1'b1;
6882: pixelout<=1'b1;
6883: pixelout<=1'b1;
6884: pixelout<=1'b1;
6885: pixelout<=1'b1;
6886: pixelout<=1'b1;
6887: pixelout<=1'b1;
6888: pixelout<=1'b1;
6889: pixelout<=1'b1;
6890: pixelout<=1'b1;
6891: pixelout<=1'b1;
6892: pixelout<=1'b1;
6893: pixelout<=1'b1;
6894: pixelout<=1'b1;
6895: pixelout<=1'b1;
6896: pixelout<=1'b1;
6897: pixelout<=1'b1;
6898: pixelout<=1'b1;
6899: pixelout<=1'b1;
6900: pixelout<=1'b1;
6901: pixelout<=1'b1;
6902: pixelout<=1'b1;
6903: pixelout<=1'b1;
6904: pixelout<=1'b1;
6905: pixelout<=1'b1;
6906: pixelout<=1'b1;
6907: pixelout<=1'b1;
6908: pixelout<=1'b1;
6909: pixelout<=1'b1;
6910: pixelout<=1'b1;
6911: pixelout<=1'b1;
6912: pixelout<=1'b1;
6913: pixelout<=1'b1;
6914: pixelout<=1'b1;
6915: pixelout<=1'b1;
6916: pixelout<=1'b1;
6917: pixelout<=1'b1;
6918: pixelout<=1'b1;
6919: pixelout<=1'b1;
6920: pixelout<=1'b1;
6921: pixelout<=1'b1;
6922: pixelout<=1'b1;
6923: pixelout<=1'b1;
6924: pixelout<=1'b1;
6925: pixelout<=1'b1;
6926: pixelout<=1'b1;
6927: pixelout<=1'b1;
6928: pixelout<=1'b1;
6929: pixelout<=1'b1;
6930: pixelout<=1'b1;
6931: pixelout<=1'b1;
6932: pixelout<=1'b1;
6933: pixelout<=1'b1;
6934: pixelout<=1'b1;
6935: pixelout<=1'b1;
6936: pixelout<=1'b1;
6937: pixelout<=1'b1;
6938: pixelout<=1'b1;
6939: pixelout<=1'b1;
6940: pixelout<=1'b1;
6941: pixelout<=1'b1;
6942: pixelout<=1'b1;
6943: pixelout<=1'b1;
6944: pixelout<=1'b1;
6945: pixelout<=1'b1;
6946: pixelout<=1'b1;
6947: pixelout<=1'b1;
6948: pixelout<=1'b1;
6949: pixelout<=1'b1;
6950: pixelout<=1'b1;
6951: pixelout<=1'b1;
6952: pixelout<=1'b1;
6953: pixelout<=1'b1;
6954: pixelout<=1'b1;
6955: pixelout<=1'b1;
6956: pixelout<=1'b1;
6957: pixelout<=1'b1;
6958: pixelout<=1'b1;
6959: pixelout<=1'b1;
6960: pixelout<=1'b1;
6961: pixelout<=1'b1;
6962: pixelout<=1'b1;
6963: pixelout<=1'b1;
6964: pixelout<=1'b1;
6965: pixelout<=1'b1;
6966: pixelout<=1'b1;
6967: pixelout<=1'b1;
6968: pixelout<=1'b1;
6969: pixelout<=1'b1;
6970: pixelout<=1'b1;
6971: pixelout<=1'b1;
6972: pixelout<=1'b1;
6973: pixelout<=1'b1;
6974: pixelout<=1'b1;
6975: pixelout<=1'b1;
6976: pixelout<=1'b1;
6977: pixelout<=1'b1;
6978: pixelout<=1'b1;
6979: pixelout<=1'b1;
6980: pixelout<=1'b1;
6981: pixelout<=1'b1;
6982: pixelout<=1'b1;
6983: pixelout<=1'b1;
6984: pixelout<=1'b1;
6985: pixelout<=1'b1;
6986: pixelout<=1'b1;
6987: pixelout<=1'b1;
6988: pixelout<=1'b1;
6989: pixelout<=1'b1;
6990: pixelout<=1'b1;
6991: pixelout<=1'b1;
6992: pixelout<=1'b1;
6993: pixelout<=1'b1;
6994: pixelout<=1'b1;
6995: pixelout<=1'b1;
6996: pixelout<=1'b1;
6997: pixelout<=1'b1;
6998: pixelout<=1'b1;
6999: pixelout<=1'b1;
7000: pixelout<=1'b1;
7001: pixelout<=1'b1;
7002: pixelout<=1'b1;
7003: pixelout<=1'b1;
7004: pixelout<=1'b1;
7005: pixelout<=1'b1;
7006: pixelout<=1'b1;
7007: pixelout<=1'b1;
7008: pixelout<=1'b1;
7009: pixelout<=1'b1;
7010: pixelout<=1'b1;
7011: pixelout<=1'b1;
7012: pixelout<=1'b1;
7013: pixelout<=1'b1;
7014: pixelout<=1'b1;
7015: pixelout<=1'b1;
7016: pixelout<=1'b1;
7017: pixelout<=1'b1;
7018: pixelout<=1'b1;
7019: pixelout<=1'b1;
7020: pixelout<=1'b1;
7021: pixelout<=1'b1;
7022: pixelout<=1'b1;
7023: pixelout<=1'b1;
7024: pixelout<=1'b1;
7025: pixelout<=1'b1;
7026: pixelout<=1'b1;
7027: pixelout<=1'b1;
7028: pixelout<=1'b1;
7029: pixelout<=1'b1;
7030: pixelout<=1'b1;
7031: pixelout<=1'b1;
7032: pixelout<=1'b1;
7033: pixelout<=1'b1;
7034: pixelout<=1'b1;
7035: pixelout<=1'b1;
7036: pixelout<=1'b1;
7037: pixelout<=1'b1;
7038: pixelout<=1'b1;
7039: pixelout<=1'b1;
7040: pixelout<=1'b1;
7041: pixelout<=1'b1;
7042: pixelout<=1'b1;
7043: pixelout<=1'b1;
7044: pixelout<=1'b1;
7045: pixelout<=1'b1;
7046: pixelout<=1'b1;
7047: pixelout<=1'b1;
7048: pixelout<=1'b1;
7049: pixelout<=1'b1;
7050: pixelout<=1'b1;
7051: pixelout<=1'b1;
7052: pixelout<=1'b1;
7053: pixelout<=1'b1;
7054: pixelout<=1'b1;
7055: pixelout<=1'b1;
7056: pixelout<=1'b1;
7057: pixelout<=1'b1;
7058: pixelout<=1'b1;
7059: pixelout<=1'b1;
7060: pixelout<=1'b1;
7061: pixelout<=1'b1;
7062: pixelout<=1'b1;
7063: pixelout<=1'b1;
7064: pixelout<=1'b1;
7065: pixelout<=1'b1;
7066: pixelout<=1'b1;
7067: pixelout<=1'b1;
7068: pixelout<=1'b1;
7069: pixelout<=1'b1;
7070: pixelout<=1'b1;
7071: pixelout<=1'b1;
7072: pixelout<=1'b1;
7073: pixelout<=1'b1;
7074: pixelout<=1'b1;
7075: pixelout<=1'b1;
7076: pixelout<=1'b1;
7077: pixelout<=1'b1;
7078: pixelout<=1'b1;
7079: pixelout<=1'b1;
7080: pixelout<=1'b1;
7081: pixelout<=1'b1;
7082: pixelout<=1'b1;
7083: pixelout<=1'b1;
7084: pixelout<=1'b1;
7085: pixelout<=1'b1;
7086: pixelout<=1'b1;
7087: pixelout<=1'b1;
7088: pixelout<=1'b1;
7089: pixelout<=1'b1;
7090: pixelout<=1'b1;
7091: pixelout<=1'b1;
7092: pixelout<=1'b1;
7093: pixelout<=1'b1;
7094: pixelout<=1'b1;
7095: pixelout<=1'b1;
7096: pixelout<=1'b1;
7097: pixelout<=1'b1;
7098: pixelout<=1'b1;
7099: pixelout<=1'b1;
7100: pixelout<=1'b1;
7101: pixelout<=1'b1;
7102: pixelout<=1'b1;
7103: pixelout<=1'b1;
7104: pixelout<=1'b1;
7105: pixelout<=1'b1;
7106: pixelout<=1'b1;
7107: pixelout<=1'b1;
7108: pixelout<=1'b1;
7109: pixelout<=1'b1;
7110: pixelout<=1'b1;
7111: pixelout<=1'b1;
7112: pixelout<=1'b1;
7113: pixelout<=1'b1;
7114: pixelout<=1'b1;
7115: pixelout<=1'b1;
7116: pixelout<=1'b1;
7117: pixelout<=1'b1;
7118: pixelout<=1'b1;
7119: pixelout<=1'b1;
7120: pixelout<=1'b1;
7121: pixelout<=1'b1;
7122: pixelout<=1'b1;
7123: pixelout<=1'b1;
7124: pixelout<=1'b1;
7125: pixelout<=1'b1;
7126: pixelout<=1'b1;
7127: pixelout<=1'b1;
7128: pixelout<=1'b1;
7129: pixelout<=1'b1;
7130: pixelout<=1'b0;
7131: pixelout<=1'b1;
7132: pixelout<=1'b1;
7133: pixelout<=1'b0;
7134: pixelout<=1'b0;
7135: pixelout<=1'b1;
7136: pixelout<=1'b1;
7137: pixelout<=1'b1;
7138: pixelout<=1'b1;
7139: pixelout<=1'b1;
7140: pixelout<=1'b1;
7141: pixelout<=1'b1;
7142: pixelout<=1'b1;
7143: pixelout<=1'b1;
7144: pixelout<=1'b1;
7145: pixelout<=1'b1;
7146: pixelout<=1'b1;
7147: pixelout<=1'b1;
7148: pixelout<=1'b1;
7149: pixelout<=1'b1;
7150: pixelout<=1'b1;
7151: pixelout<=1'b1;
7152: pixelout<=1'b1;
7153: pixelout<=1'b1;
7154: pixelout<=1'b1;
7155: pixelout<=1'b1;
7156: pixelout<=1'b1;
7157: pixelout<=1'b1;
7158: pixelout<=1'b1;
7159: pixelout<=1'b1;
7160: pixelout<=1'b1;
7161: pixelout<=1'b1;
7162: pixelout<=1'b1;
7163: pixelout<=1'b1;
7164: pixelout<=1'b1;
7165: pixelout<=1'b1;
7166: pixelout<=1'b1;
7167: pixelout<=1'b1;
7168: pixelout<=1'b1;
7169: pixelout<=1'b1;
7170: pixelout<=1'b1;
7171: pixelout<=1'b1;
7172: pixelout<=1'b1;
7173: pixelout<=1'b1;
7174: pixelout<=1'b1;
7175: pixelout<=1'b1;
7176: pixelout<=1'b1;
7177: pixelout<=1'b1;
7178: pixelout<=1'b1;
7179: pixelout<=1'b1;
7180: pixelout<=1'b1;
7181: pixelout<=1'b1;
7182: pixelout<=1'b1;
7183: pixelout<=1'b1;
7184: pixelout<=1'b1;
7185: pixelout<=1'b1;
7186: pixelout<=1'b1;
7187: pixelout<=1'b1;
7188: pixelout<=1'b1;
7189: pixelout<=1'b1;
7190: pixelout<=1'b1;
7191: pixelout<=1'b1;
7192: pixelout<=1'b1;
7193: pixelout<=1'b1;
7194: pixelout<=1'b1;
7195: pixelout<=1'b1;
7196: pixelout<=1'b1;
7197: pixelout<=1'b1;
7198: pixelout<=1'b1;
7199: pixelout<=1'b1;
7200: pixelout<=1'b1;
7201: pixelout<=1'b1;
7202: pixelout<=1'b1;
7203: pixelout<=1'b1;
7204: pixelout<=1'b1;
7205: pixelout<=1'b1;
7206: pixelout<=1'b1;
7207: pixelout<=1'b1;
7208: pixelout<=1'b1;
7209: pixelout<=1'b1;
7210: pixelout<=1'b1;
7211: pixelout<=1'b1;
7212: pixelout<=1'b1;
7213: pixelout<=1'b1;
7214: pixelout<=1'b1;
7215: pixelout<=1'b1;
7216: pixelout<=1'b1;
7217: pixelout<=1'b1;
7218: pixelout<=1'b1;
7219: pixelout<=1'b1;
7220: pixelout<=1'b1;
7221: pixelout<=1'b1;
7222: pixelout<=1'b1;
7223: pixelout<=1'b1;
7224: pixelout<=1'b1;
7225: pixelout<=1'b1;
7226: pixelout<=1'b1;
7227: pixelout<=1'b1;
7228: pixelout<=1'b1;
7229: pixelout<=1'b1;
7230: pixelout<=1'b1;
7231: pixelout<=1'b1;
7232: pixelout<=1'b1;
7233: pixelout<=1'b1;
7234: pixelout<=1'b1;
7235: pixelout<=1'b1;
7236: pixelout<=1'b1;
7237: pixelout<=1'b1;
7238: pixelout<=1'b1;
7239: pixelout<=1'b1;
7240: pixelout<=1'b1;
7241: pixelout<=1'b1;
7242: pixelout<=1'b1;
7243: pixelout<=1'b1;
7244: pixelout<=1'b1;
7245: pixelout<=1'b1;
7246: pixelout<=1'b1;
7247: pixelout<=1'b1;
7248: pixelout<=1'b1;
7249: pixelout<=1'b1;
7250: pixelout<=1'b1;
7251: pixelout<=1'b1;
7252: pixelout<=1'b1;
7253: pixelout<=1'b1;
7254: pixelout<=1'b1;
7255: pixelout<=1'b1;
7256: pixelout<=1'b1;
7257: pixelout<=1'b1;
7258: pixelout<=1'b1;
7259: pixelout<=1'b1;
7260: pixelout<=1'b1;
7261: pixelout<=1'b1;
7262: pixelout<=1'b1;
7263: pixelout<=1'b1;
7264: pixelout<=1'b1;
7265: pixelout<=1'b1;
7266: pixelout<=1'b1;
7267: pixelout<=1'b1;
7268: pixelout<=1'b1;
7269: pixelout<=1'b1;
7270: pixelout<=1'b1;
7271: pixelout<=1'b1;
7272: pixelout<=1'b1;
7273: pixelout<=1'b1;
7274: pixelout<=1'b1;
7275: pixelout<=1'b1;
7276: pixelout<=1'b1;
7277: pixelout<=1'b1;
7278: pixelout<=1'b1;
7279: pixelout<=1'b1;
7280: pixelout<=1'b1;
7281: pixelout<=1'b1;
7282: pixelout<=1'b1;
7283: pixelout<=1'b1;
7284: pixelout<=1'b1;
7285: pixelout<=1'b1;
7286: pixelout<=1'b1;
7287: pixelout<=1'b1;
7288: pixelout<=1'b1;
7289: pixelout<=1'b1;
7290: pixelout<=1'b1;
7291: pixelout<=1'b1;
7292: pixelout<=1'b1;
7293: pixelout<=1'b1;
7294: pixelout<=1'b1;
7295: pixelout<=1'b1;
7296: pixelout<=1'b1;
7297: pixelout<=1'b1;
7298: pixelout<=1'b1;
7299: pixelout<=1'b1;
7300: pixelout<=1'b1;
7301: pixelout<=1'b1;
7302: pixelout<=1'b1;
7303: pixelout<=1'b1;
7304: pixelout<=1'b1;
7305: pixelout<=1'b1;
7306: pixelout<=1'b1;
7307: pixelout<=1'b1;
7308: pixelout<=1'b1;
7309: pixelout<=1'b1;
7310: pixelout<=1'b1;
7311: pixelout<=1'b1;
7312: pixelout<=1'b1;
7313: pixelout<=1'b1;
7314: pixelout<=1'b1;
7315: pixelout<=1'b1;
7316: pixelout<=1'b1;
7317: pixelout<=1'b1;
7318: pixelout<=1'b1;
7319: pixelout<=1'b1;
7320: pixelout<=1'b1;
7321: pixelout<=1'b1;
7322: pixelout<=1'b1;
7323: pixelout<=1'b1;
7324: pixelout<=1'b1;
7325: pixelout<=1'b1;
7326: pixelout<=1'b1;
7327: pixelout<=1'b1;
7328: pixelout<=1'b1;
7329: pixelout<=1'b1;
7330: pixelout<=1'b1;
7331: pixelout<=1'b1;
7332: pixelout<=1'b1;
7333: pixelout<=1'b1;
7334: pixelout<=1'b1;
7335: pixelout<=1'b1;
7336: pixelout<=1'b1;
7337: pixelout<=1'b1;
7338: pixelout<=1'b1;
7339: pixelout<=1'b1;
7340: pixelout<=1'b1;
7341: pixelout<=1'b1;
7342: pixelout<=1'b1;
7343: pixelout<=1'b1;
7344: pixelout<=1'b1;
7345: pixelout<=1'b1;
7346: pixelout<=1'b1;
7347: pixelout<=1'b1;
7348: pixelout<=1'b1;
7349: pixelout<=1'b1;
7350: pixelout<=1'b1;
7351: pixelout<=1'b1;
7352: pixelout<=1'b1;
7353: pixelout<=1'b1;
7354: pixelout<=1'b1;
7355: pixelout<=1'b1;
7356: pixelout<=1'b1;
7357: pixelout<=1'b1;
7358: pixelout<=1'b1;
7359: pixelout<=1'b1;
7360: pixelout<=1'b1;
7361: pixelout<=1'b1;
7362: pixelout<=1'b1;
7363: pixelout<=1'b1;
7364: pixelout<=1'b1;
7365: pixelout<=1'b1;
7366: pixelout<=1'b1;
7367: pixelout<=1'b1;
7368: pixelout<=1'b1;
7369: pixelout<=1'b1;
7370: pixelout<=1'b1;
7371: pixelout<=1'b1;
7372: pixelout<=1'b1;
7373: pixelout<=1'b1;
7374: pixelout<=1'b0;
7375: pixelout<=1'b1;
7376: pixelout<=1'b1;
7377: pixelout<=1'b1;
7378: pixelout<=1'b1;
7379: pixelout<=1'b1;
7380: pixelout<=1'b1;
7381: pixelout<=1'b1;
7382: pixelout<=1'b0;
7383: pixelout<=1'b1;
7384: pixelout<=1'b1;
7385: pixelout<=1'b1;
7386: pixelout<=1'b1;
7387: pixelout<=1'b1;
7388: pixelout<=1'b1;
7389: pixelout<=1'b1;
7390: pixelout<=1'b1;
7391: pixelout<=1'b1;
7392: pixelout<=1'b1;
7393: pixelout<=1'b1;
7394: pixelout<=1'b1;
7395: pixelout<=1'b1;
7396: pixelout<=1'b1;
7397: pixelout<=1'b1;
7398: pixelout<=1'b1;
7399: pixelout<=1'b1;
7400: pixelout<=1'b1;
7401: pixelout<=1'b1;
7402: pixelout<=1'b1;
7403: pixelout<=1'b1;
7404: pixelout<=1'b1;
7405: pixelout<=1'b1;
7406: pixelout<=1'b1;
7407: pixelout<=1'b1;
7408: pixelout<=1'b1;
7409: pixelout<=1'b1;
7410: pixelout<=1'b1;
7411: pixelout<=1'b1;
7412: pixelout<=1'b1;
7413: pixelout<=1'b1;
7414: pixelout<=1'b1;
7415: pixelout<=1'b1;
7416: pixelout<=1'b1;
7417: pixelout<=1'b1;
7418: pixelout<=1'b1;
7419: pixelout<=1'b1;
7420: pixelout<=1'b1;
7421: pixelout<=1'b1;
7422: pixelout<=1'b1;
7423: pixelout<=1'b1;
7424: pixelout<=1'b1;
7425: pixelout<=1'b1;
7426: pixelout<=1'b1;
7427: pixelout<=1'b1;
7428: pixelout<=1'b1;
7429: pixelout<=1'b1;
7430: pixelout<=1'b1;
7431: pixelout<=1'b1;
7432: pixelout<=1'b1;
7433: pixelout<=1'b1;
7434: pixelout<=1'b1;
7435: pixelout<=1'b1;
7436: pixelout<=1'b1;
7437: pixelout<=1'b1;
7438: pixelout<=1'b1;
7439: pixelout<=1'b1;
7440: pixelout<=1'b1;
7441: pixelout<=1'b1;
7442: pixelout<=1'b1;
7443: pixelout<=1'b1;
7444: pixelout<=1'b1;
7445: pixelout<=1'b1;
7446: pixelout<=1'b1;
7447: pixelout<=1'b1;
7448: pixelout<=1'b1;
7449: pixelout<=1'b1;
7450: pixelout<=1'b1;
7451: pixelout<=1'b1;
7452: pixelout<=1'b1;
7453: pixelout<=1'b1;
7454: pixelout<=1'b1;
7455: pixelout<=1'b1;
7456: pixelout<=1'b1;
7457: pixelout<=1'b1;
7458: pixelout<=1'b1;
7459: pixelout<=1'b1;
7460: pixelout<=1'b1;
7461: pixelout<=1'b1;
7462: pixelout<=1'b1;
7463: pixelout<=1'b1;
7464: pixelout<=1'b1;
7465: pixelout<=1'b1;
7466: pixelout<=1'b1;
7467: pixelout<=1'b1;
7468: pixelout<=1'b1;
7469: pixelout<=1'b1;
7470: pixelout<=1'b1;
7471: pixelout<=1'b1;
7472: pixelout<=1'b1;
7473: pixelout<=1'b1;
7474: pixelout<=1'b1;
7475: pixelout<=1'b1;
7476: pixelout<=1'b1;
7477: pixelout<=1'b1;
7478: pixelout<=1'b1;
7479: pixelout<=1'b1;
7480: pixelout<=1'b1;
7481: pixelout<=1'b1;
7482: pixelout<=1'b1;
7483: pixelout<=1'b1;
7484: pixelout<=1'b1;
7485: pixelout<=1'b1;
7486: pixelout<=1'b1;
7487: pixelout<=1'b1;
7488: pixelout<=1'b1;
7489: pixelout<=1'b1;
7490: pixelout<=1'b1;
7491: pixelout<=1'b1;
7492: pixelout<=1'b1;
7493: pixelout<=1'b1;
7494: pixelout<=1'b1;
7495: pixelout<=1'b1;
7496: pixelout<=1'b1;
7497: pixelout<=1'b1;
7498: pixelout<=1'b1;
7499: pixelout<=1'b1;
7500: pixelout<=1'b1;
7501: pixelout<=1'b1;
7502: pixelout<=1'b1;
7503: pixelout<=1'b1;
7504: pixelout<=1'b1;
7505: pixelout<=1'b1;
7506: pixelout<=1'b1;
7507: pixelout<=1'b1;
7508: pixelout<=1'b1;
7509: pixelout<=1'b1;
7510: pixelout<=1'b1;
7511: pixelout<=1'b1;
7512: pixelout<=1'b1;
7513: pixelout<=1'b1;
7514: pixelout<=1'b1;
7515: pixelout<=1'b1;
7516: pixelout<=1'b1;
7517: pixelout<=1'b1;
7518: pixelout<=1'b1;
7519: pixelout<=1'b1;
7520: pixelout<=1'b1;
7521: pixelout<=1'b1;
7522: pixelout<=1'b1;
7523: pixelout<=1'b1;
7524: pixelout<=1'b1;
7525: pixelout<=1'b1;
7526: pixelout<=1'b1;
7527: pixelout<=1'b1;
7528: pixelout<=1'b1;
7529: pixelout<=1'b1;
7530: pixelout<=1'b1;
7531: pixelout<=1'b1;
7532: pixelout<=1'b1;
7533: pixelout<=1'b1;
7534: pixelout<=1'b1;
7535: pixelout<=1'b1;
7536: pixelout<=1'b1;
7537: pixelout<=1'b1;
7538: pixelout<=1'b1;
7539: pixelout<=1'b1;
7540: pixelout<=1'b1;
7541: pixelout<=1'b1;
7542: pixelout<=1'b1;
7543: pixelout<=1'b1;
7544: pixelout<=1'b1;
7545: pixelout<=1'b1;
7546: pixelout<=1'b1;
7547: pixelout<=1'b1;
7548: pixelout<=1'b1;
7549: pixelout<=1'b1;
7550: pixelout<=1'b1;
7551: pixelout<=1'b1;
7552: pixelout<=1'b1;
7553: pixelout<=1'b1;
7554: pixelout<=1'b1;
7555: pixelout<=1'b1;
7556: pixelout<=1'b1;
7557: pixelout<=1'b1;
7558: pixelout<=1'b1;
7559: pixelout<=1'b1;
7560: pixelout<=1'b1;
7561: pixelout<=1'b1;
7562: pixelout<=1'b1;
7563: pixelout<=1'b1;
7564: pixelout<=1'b1;
7565: pixelout<=1'b1;
7566: pixelout<=1'b1;
7567: pixelout<=1'b1;
7568: pixelout<=1'b1;
7569: pixelout<=1'b1;
7570: pixelout<=1'b1;
7571: pixelout<=1'b1;
7572: pixelout<=1'b1;
7573: pixelout<=1'b1;
7574: pixelout<=1'b1;
7575: pixelout<=1'b1;
7576: pixelout<=1'b1;
7577: pixelout<=1'b1;
7578: pixelout<=1'b1;
7579: pixelout<=1'b1;
7580: pixelout<=1'b1;
7581: pixelout<=1'b1;
7582: pixelout<=1'b1;
7583: pixelout<=1'b1;
7584: pixelout<=1'b1;
7585: pixelout<=1'b1;
7586: pixelout<=1'b1;
7587: pixelout<=1'b1;
7588: pixelout<=1'b1;
7589: pixelout<=1'b1;
7590: pixelout<=1'b1;
7591: pixelout<=1'b1;
7592: pixelout<=1'b1;
7593: pixelout<=1'b1;
7594: pixelout<=1'b1;
7595: pixelout<=1'b1;
7596: pixelout<=1'b1;
7597: pixelout<=1'b1;
7598: pixelout<=1'b1;
7599: pixelout<=1'b1;
7600: pixelout<=1'b1;
7601: pixelout<=1'b1;
7602: pixelout<=1'b1;
7603: pixelout<=1'b1;
7604: pixelout<=1'b1;
7605: pixelout<=1'b1;
7606: pixelout<=1'b1;
7607: pixelout<=1'b1;
7608: pixelout<=1'b1;
7609: pixelout<=1'b1;
7610: pixelout<=1'b1;
7611: pixelout<=1'b1;
7612: pixelout<=1'b1;
7613: pixelout<=1'b1;
7614: pixelout<=1'b1;
7615: pixelout<=1'b1;
7616: pixelout<=1'b1;
7617: pixelout<=1'b1;
7618: pixelout<=1'b1;
7619: pixelout<=1'b1;
7620: pixelout<=1'b1;
7621: pixelout<=1'b1;
7622: pixelout<=1'b0;
7623: pixelout<=1'b1;
7624: pixelout<=1'b1;
7625: pixelout<=1'b1;
7626: pixelout<=1'b1;
7627: pixelout<=1'b1;
7628: pixelout<=1'b1;
7629: pixelout<=1'b1;
7630: pixelout<=1'b1;
7631: pixelout<=1'b1;
7632: pixelout<=1'b1;
7633: pixelout<=1'b1;
7634: pixelout<=1'b1;
7635: pixelout<=1'b1;
7636: pixelout<=1'b1;
7637: pixelout<=1'b1;
7638: pixelout<=1'b1;
7639: pixelout<=1'b1;
7640: pixelout<=1'b1;
7641: pixelout<=1'b1;
7642: pixelout<=1'b1;
7643: pixelout<=1'b1;
7644: pixelout<=1'b1;
7645: pixelout<=1'b1;
7646: pixelout<=1'b1;
7647: pixelout<=1'b1;
7648: pixelout<=1'b1;
7649: pixelout<=1'b1;
7650: pixelout<=1'b1;
7651: pixelout<=1'b1;
7652: pixelout<=1'b1;
7653: pixelout<=1'b1;
7654: pixelout<=1'b1;
7655: pixelout<=1'b1;
7656: pixelout<=1'b1;
7657: pixelout<=1'b1;
7658: pixelout<=1'b1;
7659: pixelout<=1'b1;
7660: pixelout<=1'b1;
7661: pixelout<=1'b1;
7662: pixelout<=1'b1;
7663: pixelout<=1'b1;
7664: pixelout<=1'b1;
7665: pixelout<=1'b1;
7666: pixelout<=1'b1;
7667: pixelout<=1'b1;
7668: pixelout<=1'b1;
7669: pixelout<=1'b1;
7670: pixelout<=1'b1;
7671: pixelout<=1'b1;
7672: pixelout<=1'b1;
7673: pixelout<=1'b1;
7674: pixelout<=1'b1;
7675: pixelout<=1'b1;
7676: pixelout<=1'b1;
7677: pixelout<=1'b1;
7678: pixelout<=1'b1;
7679: pixelout<=1'b1;
7680: pixelout<=1'b1;
7681: pixelout<=1'b1;
7682: pixelout<=1'b1;
7683: pixelout<=1'b1;
7684: pixelout<=1'b1;
7685: pixelout<=1'b1;
7686: pixelout<=1'b1;
7687: pixelout<=1'b1;
7688: pixelout<=1'b1;
7689: pixelout<=1'b1;
7690: pixelout<=1'b1;
7691: pixelout<=1'b1;
7692: pixelout<=1'b1;
7693: pixelout<=1'b1;
7694: pixelout<=1'b1;
7695: pixelout<=1'b1;
7696: pixelout<=1'b1;
7697: pixelout<=1'b1;
7698: pixelout<=1'b1;
7699: pixelout<=1'b1;
7700: pixelout<=1'b1;
7701: pixelout<=1'b1;
7702: pixelout<=1'b1;
7703: pixelout<=1'b1;
7704: pixelout<=1'b1;
7705: pixelout<=1'b1;
7706: pixelout<=1'b1;
7707: pixelout<=1'b1;
7708: pixelout<=1'b1;
7709: pixelout<=1'b1;
7710: pixelout<=1'b1;
7711: pixelout<=1'b1;
7712: pixelout<=1'b1;
7713: pixelout<=1'b1;
7714: pixelout<=1'b1;
7715: pixelout<=1'b1;
7716: pixelout<=1'b1;
7717: pixelout<=1'b1;
7718: pixelout<=1'b1;
7719: pixelout<=1'b1;
7720: pixelout<=1'b1;
7721: pixelout<=1'b1;
7722: pixelout<=1'b1;
7723: pixelout<=1'b1;
7724: pixelout<=1'b1;
7725: pixelout<=1'b1;
7726: pixelout<=1'b1;
7727: pixelout<=1'b1;
7728: pixelout<=1'b1;
7729: pixelout<=1'b1;
7730: pixelout<=1'b1;
7731: pixelout<=1'b1;
7732: pixelout<=1'b1;
7733: pixelout<=1'b1;
7734: pixelout<=1'b1;
7735: pixelout<=1'b1;
7736: pixelout<=1'b1;
7737: pixelout<=1'b1;
7738: pixelout<=1'b1;
7739: pixelout<=1'b1;
7740: pixelout<=1'b1;
7741: pixelout<=1'b1;
7742: pixelout<=1'b1;
7743: pixelout<=1'b1;
7744: pixelout<=1'b1;
7745: pixelout<=1'b1;
7746: pixelout<=1'b1;
7747: pixelout<=1'b1;
7748: pixelout<=1'b1;
7749: pixelout<=1'b1;
7750: pixelout<=1'b1;
7751: pixelout<=1'b1;
7752: pixelout<=1'b1;
7753: pixelout<=1'b1;
7754: pixelout<=1'b1;
7755: pixelout<=1'b1;
7756: pixelout<=1'b1;
7757: pixelout<=1'b1;
7758: pixelout<=1'b1;
7759: pixelout<=1'b1;
7760: pixelout<=1'b1;
7761: pixelout<=1'b1;
7762: pixelout<=1'b1;
7763: pixelout<=1'b1;
7764: pixelout<=1'b1;
7765: pixelout<=1'b1;
7766: pixelout<=1'b1;
7767: pixelout<=1'b1;
7768: pixelout<=1'b1;
7769: pixelout<=1'b1;
7770: pixelout<=1'b1;
7771: pixelout<=1'b1;
7772: pixelout<=1'b1;
7773: pixelout<=1'b1;
7774: pixelout<=1'b1;
7775: pixelout<=1'b1;
7776: pixelout<=1'b1;
7777: pixelout<=1'b1;
7778: pixelout<=1'b1;
7779: pixelout<=1'b1;
7780: pixelout<=1'b1;
7781: pixelout<=1'b1;
7782: pixelout<=1'b1;
7783: pixelout<=1'b1;
7784: pixelout<=1'b1;
7785: pixelout<=1'b1;
7786: pixelout<=1'b1;
7787: pixelout<=1'b1;
7788: pixelout<=1'b1;
7789: pixelout<=1'b1;
7790: pixelout<=1'b1;
7791: pixelout<=1'b1;
7792: pixelout<=1'b1;
7793: pixelout<=1'b1;
7794: pixelout<=1'b1;
7795: pixelout<=1'b1;
7796: pixelout<=1'b1;
7797: pixelout<=1'b1;
7798: pixelout<=1'b1;
7799: pixelout<=1'b1;
7800: pixelout<=1'b1;
7801: pixelout<=1'b1;
7802: pixelout<=1'b1;
7803: pixelout<=1'b1;
7804: pixelout<=1'b1;
7805: pixelout<=1'b1;
7806: pixelout<=1'b1;
7807: pixelout<=1'b1;
7808: pixelout<=1'b1;
7809: pixelout<=1'b1;
7810: pixelout<=1'b1;
7811: pixelout<=1'b1;
7812: pixelout<=1'b1;
7813: pixelout<=1'b1;
7814: pixelout<=1'b1;
7815: pixelout<=1'b1;
7816: pixelout<=1'b1;
7817: pixelout<=1'b1;
7818: pixelout<=1'b1;
7819: pixelout<=1'b1;
7820: pixelout<=1'b1;
7821: pixelout<=1'b1;
7822: pixelout<=1'b1;
7823: pixelout<=1'b1;
7824: pixelout<=1'b1;
7825: pixelout<=1'b1;
7826: pixelout<=1'b1;
7827: pixelout<=1'b1;
7828: pixelout<=1'b1;
7829: pixelout<=1'b1;
7830: pixelout<=1'b1;
7831: pixelout<=1'b1;
7832: pixelout<=1'b1;
7833: pixelout<=1'b1;
7834: pixelout<=1'b1;
7835: pixelout<=1'b1;
7836: pixelout<=1'b1;
7837: pixelout<=1'b1;
7838: pixelout<=1'b1;
7839: pixelout<=1'b1;
7840: pixelout<=1'b1;
7841: pixelout<=1'b1;
7842: pixelout<=1'b1;
7843: pixelout<=1'b1;
7844: pixelout<=1'b1;
7845: pixelout<=1'b1;
7846: pixelout<=1'b1;
7847: pixelout<=1'b1;
7848: pixelout<=1'b1;
7849: pixelout<=1'b1;
7850: pixelout<=1'b1;
7851: pixelout<=1'b1;
7852: pixelout<=1'b1;
7853: pixelout<=1'b1;
7854: pixelout<=1'b1;
7855: pixelout<=1'b1;
7856: pixelout<=1'b1;
7857: pixelout<=1'b1;
7858: pixelout<=1'b1;
7859: pixelout<=1'b1;
7860: pixelout<=1'b1;
7861: pixelout<=1'b1;
7862: pixelout<=1'b0;
7863: pixelout<=1'b1;
7864: pixelout<=1'b1;
7865: pixelout<=1'b1;
7866: pixelout<=1'b1;
7867: pixelout<=1'b1;
7868: pixelout<=1'b1;
7869: pixelout<=1'b1;
7870: pixelout<=1'b1;
7871: pixelout<=1'b1;
7872: pixelout<=1'b1;
7873: pixelout<=1'b1;
7874: pixelout<=1'b1;
7875: pixelout<=1'b1;
7876: pixelout<=1'b1;
7877: pixelout<=1'b1;
7878: pixelout<=1'b1;
7879: pixelout<=1'b1;
7880: pixelout<=1'b1;
7881: pixelout<=1'b1;
7882: pixelout<=1'b1;
7883: pixelout<=1'b1;
7884: pixelout<=1'b1;
7885: pixelout<=1'b1;
7886: pixelout<=1'b1;
7887: pixelout<=1'b1;
7888: pixelout<=1'b1;
7889: pixelout<=1'b1;
7890: pixelout<=1'b1;
7891: pixelout<=1'b1;
7892: pixelout<=1'b1;
7893: pixelout<=1'b1;
7894: pixelout<=1'b1;
7895: pixelout<=1'b1;
7896: pixelout<=1'b1;
7897: pixelout<=1'b1;
7898: pixelout<=1'b1;
7899: pixelout<=1'b1;
7900: pixelout<=1'b1;
7901: pixelout<=1'b1;
7902: pixelout<=1'b1;
7903: pixelout<=1'b1;
7904: pixelout<=1'b1;
7905: pixelout<=1'b1;
7906: pixelout<=1'b1;
7907: pixelout<=1'b1;
7908: pixelout<=1'b1;
7909: pixelout<=1'b1;
7910: pixelout<=1'b1;
7911: pixelout<=1'b1;
7912: pixelout<=1'b1;
7913: pixelout<=1'b1;
7914: pixelout<=1'b1;
7915: pixelout<=1'b1;
7916: pixelout<=1'b1;
7917: pixelout<=1'b1;
7918: pixelout<=1'b1;
7919: pixelout<=1'b1;
7920: pixelout<=1'b1;
7921: pixelout<=1'b1;
7922: pixelout<=1'b1;
7923: pixelout<=1'b1;
7924: pixelout<=1'b1;
7925: pixelout<=1'b1;
7926: pixelout<=1'b1;
7927: pixelout<=1'b1;
7928: pixelout<=1'b1;
7929: pixelout<=1'b1;
7930: pixelout<=1'b1;
7931: pixelout<=1'b1;
7932: pixelout<=1'b1;
7933: pixelout<=1'b1;
7934: pixelout<=1'b1;
7935: pixelout<=1'b1;
7936: pixelout<=1'b1;
7937: pixelout<=1'b1;
7938: pixelout<=1'b1;
7939: pixelout<=1'b1;
7940: pixelout<=1'b1;
7941: pixelout<=1'b1;
7942: pixelout<=1'b1;
7943: pixelout<=1'b1;
7944: pixelout<=1'b1;
7945: pixelout<=1'b1;
7946: pixelout<=1'b1;
7947: pixelout<=1'b1;
7948: pixelout<=1'b1;
7949: pixelout<=1'b1;
7950: pixelout<=1'b1;
7951: pixelout<=1'b1;
7952: pixelout<=1'b1;
7953: pixelout<=1'b1;
7954: pixelout<=1'b1;
7955: pixelout<=1'b1;
7956: pixelout<=1'b1;
7957: pixelout<=1'b1;
7958: pixelout<=1'b1;
7959: pixelout<=1'b1;
7960: pixelout<=1'b1;
7961: pixelout<=1'b1;
7962: pixelout<=1'b1;
7963: pixelout<=1'b1;
7964: pixelout<=1'b1;
7965: pixelout<=1'b1;
7966: pixelout<=1'b1;
7967: pixelout<=1'b1;
7968: pixelout<=1'b1;
7969: pixelout<=1'b1;
7970: pixelout<=1'b1;
7971: pixelout<=1'b1;
7972: pixelout<=1'b1;
7973: pixelout<=1'b1;
7974: pixelout<=1'b1;
7975: pixelout<=1'b1;
7976: pixelout<=1'b1;
7977: pixelout<=1'b1;
7978: pixelout<=1'b1;
7979: pixelout<=1'b1;
7980: pixelout<=1'b1;
7981: pixelout<=1'b1;
7982: pixelout<=1'b1;
7983: pixelout<=1'b1;
7984: pixelout<=1'b1;
7985: pixelout<=1'b1;
7986: pixelout<=1'b1;
7987: pixelout<=1'b1;
7988: pixelout<=1'b1;
7989: pixelout<=1'b1;
7990: pixelout<=1'b1;
7991: pixelout<=1'b1;
7992: pixelout<=1'b0;
7993: pixelout<=1'b1;
7994: pixelout<=1'b1;
7995: pixelout<=1'b1;
7996: pixelout<=1'b1;
7997: pixelout<=1'b1;
7998: pixelout<=1'b1;
7999: pixelout<=1'b1;
8000: pixelout<=1'b1;
8001: pixelout<=1'b1;
8002: pixelout<=1'b1;
8003: pixelout<=1'b1;
8004: pixelout<=1'b1;
8005: pixelout<=1'b1;
8006: pixelout<=1'b1;
8007: pixelout<=1'b1;
8008: pixelout<=1'b1;
8009: pixelout<=1'b1;
8010: pixelout<=1'b1;
8011: pixelout<=1'b1;
8012: pixelout<=1'b1;
8013: pixelout<=1'b1;
8014: pixelout<=1'b1;
8015: pixelout<=1'b1;
8016: pixelout<=1'b1;
8017: pixelout<=1'b1;
8018: pixelout<=1'b1;
8019: pixelout<=1'b1;
8020: pixelout<=1'b1;
8021: pixelout<=1'b1;
8022: pixelout<=1'b0;
8023: pixelout<=1'b0;
8024: pixelout<=1'b0;
8025: pixelout<=1'b0;
8026: pixelout<=1'b0;
8027: pixelout<=1'b1;
8028: pixelout<=1'b0;
8029: pixelout<=1'b1;
8030: pixelout<=1'b1;
8031: pixelout<=1'b1;
8032: pixelout<=1'b1;
8033: pixelout<=1'b1;
8034: pixelout<=1'b1;
8035: pixelout<=1'b1;
8036: pixelout<=1'b1;
8037: pixelout<=1'b1;
8038: pixelout<=1'b1;
8039: pixelout<=1'b1;
8040: pixelout<=1'b1;
8041: pixelout<=1'b1;
8042: pixelout<=1'b0;
8043: pixelout<=1'b1;
8044: pixelout<=1'b1;
8045: pixelout<=1'b1;
8046: pixelout<=1'b1;
8047: pixelout<=1'b0;
8048: pixelout<=1'b0;
8049: pixelout<=1'b0;
8050: pixelout<=1'b0;
8051: pixelout<=1'b1;
8052: pixelout<=1'b1;
8053: pixelout<=1'b1;
8054: pixelout<=1'b1;
8055: pixelout<=1'b1;
8056: pixelout<=1'b1;
8057: pixelout<=1'b1;
8058: pixelout<=1'b1;
8059: pixelout<=1'b1;
8060: pixelout<=1'b1;
8061: pixelout<=1'b1;
8062: pixelout<=1'b1;
8063: pixelout<=1'b1;
8064: pixelout<=1'b1;
8065: pixelout<=1'b1;
8066: pixelout<=1'b1;
8067: pixelout<=1'b1;
8068: pixelout<=1'b1;
8069: pixelout<=1'b1;
8070: pixelout<=1'b1;
8071: pixelout<=1'b1;
8072: pixelout<=1'b1;
8073: pixelout<=1'b1;
8074: pixelout<=1'b1;
8075: pixelout<=1'b1;
8076: pixelout<=1'b1;
8077: pixelout<=1'b1;
8078: pixelout<=1'b1;
8079: pixelout<=1'b1;
8080: pixelout<=1'b1;
8081: pixelout<=1'b1;
8082: pixelout<=1'b1;
8083: pixelout<=1'b1;
8084: pixelout<=1'b1;
8085: pixelout<=1'b1;
8086: pixelout<=1'b1;
8087: pixelout<=1'b1;
8088: pixelout<=1'b1;
8089: pixelout<=1'b1;
8090: pixelout<=1'b1;
8091: pixelout<=1'b1;
8092: pixelout<=1'b1;
8093: pixelout<=1'b1;
8094: pixelout<=1'b1;
8095: pixelout<=1'b1;
8096: pixelout<=1'b1;
8097: pixelout<=1'b1;
8098: pixelout<=1'b1;
8099: pixelout<=1'b1;
8100: pixelout<=1'b1;
8101: pixelout<=1'b1;
8102: pixelout<=1'b0;
8103: pixelout<=1'b1;
8104: pixelout<=1'b1;
8105: pixelout<=1'b1;
8106: pixelout<=1'b1;
8107: pixelout<=1'b1;
8108: pixelout<=1'b1;
8109: pixelout<=1'b1;
8110: pixelout<=1'b1;
8111: pixelout<=1'b1;
8112: pixelout<=1'b1;
8113: pixelout<=1'b1;
8114: pixelout<=1'b1;
8115: pixelout<=1'b1;
8116: pixelout<=1'b1;
8117: pixelout<=1'b1;
8118: pixelout<=1'b1;
8119: pixelout<=1'b1;
8120: pixelout<=1'b1;
8121: pixelout<=1'b1;
8122: pixelout<=1'b1;
8123: pixelout<=1'b1;
8124: pixelout<=1'b1;
8125: pixelout<=1'b1;
8126: pixelout<=1'b1;
8127: pixelout<=1'b1;
8128: pixelout<=1'b1;
8129: pixelout<=1'b1;
8130: pixelout<=1'b1;
8131: pixelout<=1'b1;
8132: pixelout<=1'b1;
8133: pixelout<=1'b1;
8134: pixelout<=1'b1;
8135: pixelout<=1'b1;
8136: pixelout<=1'b1;
8137: pixelout<=1'b1;
8138: pixelout<=1'b1;
8139: pixelout<=1'b1;
8140: pixelout<=1'b1;
8141: pixelout<=1'b1;
8142: pixelout<=1'b1;
8143: pixelout<=1'b1;
8144: pixelout<=1'b1;
8145: pixelout<=1'b1;
8146: pixelout<=1'b1;
8147: pixelout<=1'b1;
8148: pixelout<=1'b1;
8149: pixelout<=1'b1;
8150: pixelout<=1'b1;
8151: pixelout<=1'b1;
8152: pixelout<=1'b1;
8153: pixelout<=1'b1;
8154: pixelout<=1'b1;
8155: pixelout<=1'b1;
8156: pixelout<=1'b1;
8157: pixelout<=1'b1;
8158: pixelout<=1'b1;
8159: pixelout<=1'b1;
8160: pixelout<=1'b1;
8161: pixelout<=1'b1;
8162: pixelout<=1'b1;
8163: pixelout<=1'b1;
8164: pixelout<=1'b1;
8165: pixelout<=1'b1;
8166: pixelout<=1'b1;
8167: pixelout<=1'b1;
8168: pixelout<=1'b1;
8169: pixelout<=1'b1;
8170: pixelout<=1'b1;
8171: pixelout<=1'b1;
8172: pixelout<=1'b1;
8173: pixelout<=1'b1;
8174: pixelout<=1'b1;
8175: pixelout<=1'b1;
8176: pixelout<=1'b1;
8177: pixelout<=1'b1;
8178: pixelout<=1'b1;
8179: pixelout<=1'b1;
8180: pixelout<=1'b1;
8181: pixelout<=1'b1;
8182: pixelout<=1'b1;
8183: pixelout<=1'b1;
8184: pixelout<=1'b1;
8185: pixelout<=1'b1;
8186: pixelout<=1'b1;
8187: pixelout<=1'b1;
8188: pixelout<=1'b1;
8189: pixelout<=1'b1;
8190: pixelout<=1'b1;
8191: pixelout<=1'b1;
8192: pixelout<=1'b1;
8193: pixelout<=1'b1;
8194: pixelout<=1'b1;
8195: pixelout<=1'b1;
8196: pixelout<=1'b1;
8197: pixelout<=1'b1;
8198: pixelout<=1'b1;
8199: pixelout<=1'b1;
8200: pixelout<=1'b1;
8201: pixelout<=1'b1;
8202: pixelout<=1'b1;
8203: pixelout<=1'b1;
8204: pixelout<=1'b1;
8205: pixelout<=1'b1;
8206: pixelout<=1'b1;
8207: pixelout<=1'b1;
8208: pixelout<=1'b1;
8209: pixelout<=1'b1;
8210: pixelout<=1'b1;
8211: pixelout<=1'b1;
8212: pixelout<=1'b1;
8213: pixelout<=1'b1;
8214: pixelout<=1'b1;
8215: pixelout<=1'b1;
8216: pixelout<=1'b1;
8217: pixelout<=1'b1;
8218: pixelout<=1'b1;
8219: pixelout<=1'b1;
8220: pixelout<=1'b1;
8221: pixelout<=1'b1;
8222: pixelout<=1'b1;
8223: pixelout<=1'b1;
8224: pixelout<=1'b1;
8225: pixelout<=1'b1;
8226: pixelout<=1'b1;
8227: pixelout<=1'b1;
8228: pixelout<=1'b1;
8229: pixelout<=1'b1;
8230: pixelout<=1'b1;
8231: pixelout<=1'b1;
8232: pixelout<=1'b0;
8233: pixelout<=1'b1;
8234: pixelout<=1'b1;
8235: pixelout<=1'b1;
8236: pixelout<=1'b1;
8237: pixelout<=1'b1;
8238: pixelout<=1'b1;
8239: pixelout<=1'b1;
8240: pixelout<=1'b1;
8241: pixelout<=1'b1;
8242: pixelout<=1'b1;
8243: pixelout<=1'b1;
8244: pixelout<=1'b1;
8245: pixelout<=1'b1;
8246: pixelout<=1'b1;
8247: pixelout<=1'b1;
8248: pixelout<=1'b1;
8249: pixelout<=1'b1;
8250: pixelout<=1'b1;
8251: pixelout<=1'b1;
8252: pixelout<=1'b1;
8253: pixelout<=1'b1;
8254: pixelout<=1'b1;
8255: pixelout<=1'b1;
8256: pixelout<=1'b1;
8257: pixelout<=1'b1;
8258: pixelout<=1'b1;
8259: pixelout<=1'b1;
8260: pixelout<=1'b1;
8261: pixelout<=1'b1;
8262: pixelout<=1'b0;
8263: pixelout<=1'b1;
8264: pixelout<=1'b1;
8265: pixelout<=1'b1;
8266: pixelout<=1'b1;
8267: pixelout<=1'b1;
8268: pixelout<=1'b1;
8269: pixelout<=1'b1;
8270: pixelout<=1'b1;
8271: pixelout<=1'b1;
8272: pixelout<=1'b1;
8273: pixelout<=1'b1;
8274: pixelout<=1'b1;
8275: pixelout<=1'b1;
8276: pixelout<=1'b1;
8277: pixelout<=1'b1;
8278: pixelout<=1'b1;
8279: pixelout<=1'b1;
8280: pixelout<=1'b1;
8281: pixelout<=1'b1;
8282: pixelout<=1'b1;
8283: pixelout<=1'b1;
8284: pixelout<=1'b1;
8285: pixelout<=1'b1;
8286: pixelout<=1'b1;
8287: pixelout<=1'b0;
8288: pixelout<=1'b1;
8289: pixelout<=1'b1;
8290: pixelout<=1'b1;
8291: pixelout<=1'b0;
8292: pixelout<=1'b1;
8293: pixelout<=1'b1;
8294: pixelout<=1'b1;
8295: pixelout<=1'b1;
8296: pixelout<=1'b1;
8297: pixelout<=1'b1;
8298: pixelout<=1'b1;
8299: pixelout<=1'b1;
8300: pixelout<=1'b1;
8301: pixelout<=1'b1;
8302: pixelout<=1'b1;
8303: pixelout<=1'b1;
8304: pixelout<=1'b1;
8305: pixelout<=1'b1;
8306: pixelout<=1'b1;
8307: pixelout<=1'b1;
8308: pixelout<=1'b1;
8309: pixelout<=1'b1;
8310: pixelout<=1'b1;
8311: pixelout<=1'b1;
8312: pixelout<=1'b1;
8313: pixelout<=1'b1;
8314: pixelout<=1'b1;
8315: pixelout<=1'b1;
8316: pixelout<=1'b1;
8317: pixelout<=1'b1;
8318: pixelout<=1'b1;
8319: pixelout<=1'b1;
8320: pixelout<=1'b1;
8321: pixelout<=1'b1;
8322: pixelout<=1'b1;
8323: pixelout<=1'b0;
8324: pixelout<=1'b1;
8325: pixelout<=1'b1;
8326: pixelout<=1'b1;
8327: pixelout<=1'b1;
8328: pixelout<=1'b1;
8329: pixelout<=1'b1;
8330: pixelout<=1'b1;
8331: pixelout<=1'b1;
8332: pixelout<=1'b1;
8333: pixelout<=1'b1;
8334: pixelout<=1'b1;
8335: pixelout<=1'b1;
8336: pixelout<=1'b1;
8337: pixelout<=1'b1;
8338: pixelout<=1'b0;
8339: pixelout<=1'b0;
8340: pixelout<=1'b1;
8341: pixelout<=1'b1;
8342: pixelout<=1'b0;
8343: pixelout<=1'b1;
8344: pixelout<=1'b1;
8345: pixelout<=1'b1;
8346: pixelout<=1'b1;
8347: pixelout<=1'b1;
8348: pixelout<=1'b1;
8349: pixelout<=1'b1;
8350: pixelout<=1'b1;
8351: pixelout<=1'b1;
8352: pixelout<=1'b1;
8353: pixelout<=1'b1;
8354: pixelout<=1'b1;
8355: pixelout<=1'b1;
8356: pixelout<=1'b1;
8357: pixelout<=1'b1;
8358: pixelout<=1'b1;
8359: pixelout<=1'b1;
8360: pixelout<=1'b1;
8361: pixelout<=1'b1;
8362: pixelout<=1'b1;
8363: pixelout<=1'b1;
8364: pixelout<=1'b1;
8365: pixelout<=1'b1;
8366: pixelout<=1'b1;
8367: pixelout<=1'b1;
8368: pixelout<=1'b1;
8369: pixelout<=1'b1;
8370: pixelout<=1'b1;
8371: pixelout<=1'b1;
8372: pixelout<=1'b1;
8373: pixelout<=1'b1;
8374: pixelout<=1'b1;
8375: pixelout<=1'b1;
8376: pixelout<=1'b1;
8377: pixelout<=1'b1;
8378: pixelout<=1'b1;
8379: pixelout<=1'b1;
8380: pixelout<=1'b1;
8381: pixelout<=1'b1;
8382: pixelout<=1'b1;
8383: pixelout<=1'b1;
8384: pixelout<=1'b1;
8385: pixelout<=1'b1;
8386: pixelout<=1'b1;
8387: pixelout<=1'b1;
8388: pixelout<=1'b1;
8389: pixelout<=1'b1;
8390: pixelout<=1'b1;
8391: pixelout<=1'b1;
8392: pixelout<=1'b1;
8393: pixelout<=1'b1;
8394: pixelout<=1'b1;
8395: pixelout<=1'b1;
8396: pixelout<=1'b1;
8397: pixelout<=1'b1;
8398: pixelout<=1'b1;
8399: pixelout<=1'b1;
8400: pixelout<=1'b1;
8401: pixelout<=1'b1;
8402: pixelout<=1'b1;
8403: pixelout<=1'b1;
8404: pixelout<=1'b1;
8405: pixelout<=1'b1;
8406: pixelout<=1'b1;
8407: pixelout<=1'b1;
8408: pixelout<=1'b1;
8409: pixelout<=1'b1;
8410: pixelout<=1'b1;
8411: pixelout<=1'b1;
8412: pixelout<=1'b1;
8413: pixelout<=1'b1;
8414: pixelout<=1'b1;
8415: pixelout<=1'b1;
8416: pixelout<=1'b1;
8417: pixelout<=1'b1;
8418: pixelout<=1'b1;
8419: pixelout<=1'b1;
8420: pixelout<=1'b1;
8421: pixelout<=1'b1;
8422: pixelout<=1'b1;
8423: pixelout<=1'b1;
8424: pixelout<=1'b1;
8425: pixelout<=1'b1;
8426: pixelout<=1'b1;
8427: pixelout<=1'b1;
8428: pixelout<=1'b1;
8429: pixelout<=1'b1;
8430: pixelout<=1'b1;
8431: pixelout<=1'b1;
8432: pixelout<=1'b1;
8433: pixelout<=1'b1;
8434: pixelout<=1'b1;
8435: pixelout<=1'b1;
8436: pixelout<=1'b1;
8437: pixelout<=1'b1;
8438: pixelout<=1'b1;
8439: pixelout<=1'b1;
8440: pixelout<=1'b1;
8441: pixelout<=1'b1;
8442: pixelout<=1'b1;
8443: pixelout<=1'b1;
8444: pixelout<=1'b1;
8445: pixelout<=1'b1;
8446: pixelout<=1'b1;
8447: pixelout<=1'b1;
8448: pixelout<=1'b1;
8449: pixelout<=1'b1;
8450: pixelout<=1'b1;
8451: pixelout<=1'b1;
8452: pixelout<=1'b1;
8453: pixelout<=1'b1;
8454: pixelout<=1'b1;
8455: pixelout<=1'b1;
8456: pixelout<=1'b1;
8457: pixelout<=1'b1;
8458: pixelout<=1'b1;
8459: pixelout<=1'b1;
8460: pixelout<=1'b1;
8461: pixelout<=1'b1;
8462: pixelout<=1'b1;
8463: pixelout<=1'b1;
8464: pixelout<=1'b1;
8465: pixelout<=1'b1;
8466: pixelout<=1'b1;
8467: pixelout<=1'b1;
8468: pixelout<=1'b1;
8469: pixelout<=1'b1;
8470: pixelout<=1'b1;
8471: pixelout<=1'b1;
8472: pixelout<=1'b0;
8473: pixelout<=1'b1;
8474: pixelout<=1'b1;
8475: pixelout<=1'b1;
8476: pixelout<=1'b1;
8477: pixelout<=1'b1;
8478: pixelout<=1'b1;
8479: pixelout<=1'b1;
8480: pixelout<=1'b1;
8481: pixelout<=1'b1;
8482: pixelout<=1'b1;
8483: pixelout<=1'b1;
8484: pixelout<=1'b1;
8485: pixelout<=1'b1;
8486: pixelout<=1'b1;
8487: pixelout<=1'b1;
8488: pixelout<=1'b1;
8489: pixelout<=1'b1;
8490: pixelout<=1'b1;
8491: pixelout<=1'b1;
8492: pixelout<=1'b1;
8493: pixelout<=1'b1;
8494: pixelout<=1'b1;
8495: pixelout<=1'b1;
8496: pixelout<=1'b1;
8497: pixelout<=1'b1;
8498: pixelout<=1'b1;
8499: pixelout<=1'b1;
8500: pixelout<=1'b1;
8501: pixelout<=1'b1;
8502: pixelout<=1'b0;
8503: pixelout<=1'b1;
8504: pixelout<=1'b1;
8505: pixelout<=1'b1;
8506: pixelout<=1'b1;
8507: pixelout<=1'b1;
8508: pixelout<=1'b1;
8509: pixelout<=1'b1;
8510: pixelout<=1'b1;
8511: pixelout<=1'b1;
8512: pixelout<=1'b1;
8513: pixelout<=1'b1;
8514: pixelout<=1'b1;
8515: pixelout<=1'b1;
8516: pixelout<=1'b1;
8517: pixelout<=1'b1;
8518: pixelout<=1'b1;
8519: pixelout<=1'b1;
8520: pixelout<=1'b1;
8521: pixelout<=1'b1;
8522: pixelout<=1'b1;
8523: pixelout<=1'b1;
8524: pixelout<=1'b1;
8525: pixelout<=1'b1;
8526: pixelout<=1'b1;
8527: pixelout<=1'b0;
8528: pixelout<=1'b1;
8529: pixelout<=1'b1;
8530: pixelout<=1'b1;
8531: pixelout<=1'b0;
8532: pixelout<=1'b1;
8533: pixelout<=1'b1;
8534: pixelout<=1'b1;
8535: pixelout<=1'b1;
8536: pixelout<=1'b1;
8537: pixelout<=1'b1;
8538: pixelout<=1'b1;
8539: pixelout<=1'b1;
8540: pixelout<=1'b1;
8541: pixelout<=1'b1;
8542: pixelout<=1'b1;
8543: pixelout<=1'b1;
8544: pixelout<=1'b1;
8545: pixelout<=1'b1;
8546: pixelout<=1'b1;
8547: pixelout<=1'b1;
8548: pixelout<=1'b1;
8549: pixelout<=1'b1;
8550: pixelout<=1'b1;
8551: pixelout<=1'b1;
8552: pixelout<=1'b1;
8553: pixelout<=1'b1;
8554: pixelout<=1'b1;
8555: pixelout<=1'b1;
8556: pixelout<=1'b1;
8557: pixelout<=1'b1;
8558: pixelout<=1'b1;
8559: pixelout<=1'b1;
8560: pixelout<=1'b1;
8561: pixelout<=1'b1;
8562: pixelout<=1'b1;
8563: pixelout<=1'b0;
8564: pixelout<=1'b1;
8565: pixelout<=1'b1;
8566: pixelout<=1'b1;
8567: pixelout<=1'b1;
8568: pixelout<=1'b1;
8569: pixelout<=1'b1;
8570: pixelout<=1'b1;
8571: pixelout<=1'b1;
8572: pixelout<=1'b1;
8573: pixelout<=1'b1;
8574: pixelout<=1'b1;
8575: pixelout<=1'b1;
8576: pixelout<=1'b1;
8577: pixelout<=1'b1;
8578: pixelout<=1'b0;
8579: pixelout<=1'b1;
8580: pixelout<=1'b1;
8581: pixelout<=1'b1;
8582: pixelout<=1'b0;
8583: pixelout<=1'b1;
8584: pixelout<=1'b1;
8585: pixelout<=1'b1;
8586: pixelout<=1'b1;
8587: pixelout<=1'b1;
8588: pixelout<=1'b1;
8589: pixelout<=1'b1;
8590: pixelout<=1'b1;
8591: pixelout<=1'b1;
8592: pixelout<=1'b1;
8593: pixelout<=1'b1;
8594: pixelout<=1'b1;
8595: pixelout<=1'b1;
8596: pixelout<=1'b1;
8597: pixelout<=1'b1;
8598: pixelout<=1'b1;
8599: pixelout<=1'b1;
8600: pixelout<=1'b1;
8601: pixelout<=1'b1;
8602: pixelout<=1'b1;
8603: pixelout<=1'b1;
8604: pixelout<=1'b1;
8605: pixelout<=1'b1;
8606: pixelout<=1'b1;
8607: pixelout<=1'b1;
8608: pixelout<=1'b1;
8609: pixelout<=1'b1;
8610: pixelout<=1'b1;
8611: pixelout<=1'b1;
8612: pixelout<=1'b1;
8613: pixelout<=1'b1;
8614: pixelout<=1'b1;
8615: pixelout<=1'b1;
8616: pixelout<=1'b1;
8617: pixelout<=1'b1;
8618: pixelout<=1'b1;
8619: pixelout<=1'b1;
8620: pixelout<=1'b1;
8621: pixelout<=1'b1;
8622: pixelout<=1'b1;
8623: pixelout<=1'b1;
8624: pixelout<=1'b1;
8625: pixelout<=1'b1;
8626: pixelout<=1'b1;
8627: pixelout<=1'b1;
8628: pixelout<=1'b1;
8629: pixelout<=1'b1;
8630: pixelout<=1'b1;
8631: pixelout<=1'b1;
8632: pixelout<=1'b1;
8633: pixelout<=1'b1;
8634: pixelout<=1'b1;
8635: pixelout<=1'b1;
8636: pixelout<=1'b1;
8637: pixelout<=1'b1;
8638: pixelout<=1'b1;
8639: pixelout<=1'b1;
8640: pixelout<=1'b1;
8641: pixelout<=1'b1;
8642: pixelout<=1'b1;
8643: pixelout<=1'b1;
8644: pixelout<=1'b1;
8645: pixelout<=1'b1;
8646: pixelout<=1'b1;
8647: pixelout<=1'b1;
8648: pixelout<=1'b1;
8649: pixelout<=1'b1;
8650: pixelout<=1'b1;
8651: pixelout<=1'b1;
8652: pixelout<=1'b1;
8653: pixelout<=1'b1;
8654: pixelout<=1'b1;
8655: pixelout<=1'b1;
8656: pixelout<=1'b1;
8657: pixelout<=1'b1;
8658: pixelout<=1'b1;
8659: pixelout<=1'b1;
8660: pixelout<=1'b1;
8661: pixelout<=1'b1;
8662: pixelout<=1'b1;
8663: pixelout<=1'b1;
8664: pixelout<=1'b1;
8665: pixelout<=1'b1;
8666: pixelout<=1'b1;
8667: pixelout<=1'b1;
8668: pixelout<=1'b1;
8669: pixelout<=1'b1;
8670: pixelout<=1'b1;
8671: pixelout<=1'b1;
8672: pixelout<=1'b1;
8673: pixelout<=1'b1;
8674: pixelout<=1'b1;
8675: pixelout<=1'b1;
8676: pixelout<=1'b1;
8677: pixelout<=1'b1;
8678: pixelout<=1'b1;
8679: pixelout<=1'b1;
8680: pixelout<=1'b1;
8681: pixelout<=1'b1;
8682: pixelout<=1'b1;
8683: pixelout<=1'b1;
8684: pixelout<=1'b1;
8685: pixelout<=1'b1;
8686: pixelout<=1'b1;
8687: pixelout<=1'b1;
8688: pixelout<=1'b1;
8689: pixelout<=1'b1;
8690: pixelout<=1'b1;
8691: pixelout<=1'b1;
8692: pixelout<=1'b1;
8693: pixelout<=1'b1;
8694: pixelout<=1'b1;
8695: pixelout<=1'b1;
8696: pixelout<=1'b1;
8697: pixelout<=1'b0;
8698: pixelout<=1'b0;
8699: pixelout<=1'b0;
8700: pixelout<=1'b0;
8701: pixelout<=1'b1;
8702: pixelout<=1'b0;
8703: pixelout<=1'b0;
8704: pixelout<=1'b0;
8705: pixelout<=1'b1;
8706: pixelout<=1'b1;
8707: pixelout<=1'b1;
8708: pixelout<=1'b1;
8709: pixelout<=1'b0;
8710: pixelout<=1'b0;
8711: pixelout<=1'b0;
8712: pixelout<=1'b0;
8713: pixelout<=1'b1;
8714: pixelout<=1'b1;
8715: pixelout<=1'b1;
8716: pixelout<=1'b0;
8717: pixelout<=1'b1;
8718: pixelout<=1'b1;
8719: pixelout<=1'b1;
8720: pixelout<=1'b0;
8721: pixelout<=1'b1;
8722: pixelout<=1'b1;
8723: pixelout<=1'b0;
8724: pixelout<=1'b0;
8725: pixelout<=1'b0;
8726: pixelout<=1'b1;
8727: pixelout<=1'b1;
8728: pixelout<=1'b0;
8729: pixelout<=1'b1;
8730: pixelout<=1'b1;
8731: pixelout<=1'b0;
8732: pixelout<=1'b1;
8733: pixelout<=1'b1;
8734: pixelout<=1'b1;
8735: pixelout<=1'b1;
8736: pixelout<=1'b1;
8737: pixelout<=1'b0;
8738: pixelout<=1'b1;
8739: pixelout<=1'b1;
8740: pixelout<=1'b1;
8741: pixelout<=1'b1;
8742: pixelout<=1'b0;
8743: pixelout<=1'b0;
8744: pixelout<=1'b0;
8745: pixelout<=1'b0;
8746: pixelout<=1'b1;
8747: pixelout<=1'b1;
8748: pixelout<=1'b0;
8749: pixelout<=1'b1;
8750: pixelout<=1'b0;
8751: pixelout<=1'b0;
8752: pixelout<=1'b0;
8753: pixelout<=1'b1;
8754: pixelout<=1'b1;
8755: pixelout<=1'b1;
8756: pixelout<=1'b1;
8757: pixelout<=1'b0;
8758: pixelout<=1'b0;
8759: pixelout<=1'b0;
8760: pixelout<=1'b1;
8761: pixelout<=1'b1;
8762: pixelout<=1'b1;
8763: pixelout<=1'b1;
8764: pixelout<=1'b1;
8765: pixelout<=1'b1;
8766: pixelout<=1'b1;
8767: pixelout<=1'b0;
8768: pixelout<=1'b1;
8769: pixelout<=1'b1;
8770: pixelout<=1'b1;
8771: pixelout<=1'b0;
8772: pixelout<=1'b1;
8773: pixelout<=1'b0;
8774: pixelout<=1'b1;
8775: pixelout<=1'b0;
8776: pixelout<=1'b0;
8777: pixelout<=1'b1;
8778: pixelout<=1'b1;
8779: pixelout<=1'b1;
8780: pixelout<=1'b0;
8781: pixelout<=1'b0;
8782: pixelout<=1'b1;
8783: pixelout<=1'b1;
8784: pixelout<=1'b1;
8785: pixelout<=1'b1;
8786: pixelout<=1'b1;
8787: pixelout<=1'b1;
8788: pixelout<=1'b0;
8789: pixelout<=1'b1;
8790: pixelout<=1'b1;
8791: pixelout<=1'b0;
8792: pixelout<=1'b0;
8793: pixelout<=1'b0;
8794: pixelout<=1'b1;
8795: pixelout<=1'b1;
8796: pixelout<=1'b1;
8797: pixelout<=1'b0;
8798: pixelout<=1'b0;
8799: pixelout<=1'b0;
8800: pixelout<=1'b1;
8801: pixelout<=1'b1;
8802: pixelout<=1'b1;
8803: pixelout<=1'b0;
8804: pixelout<=1'b0;
8805: pixelout<=1'b0;
8806: pixelout<=1'b1;
8807: pixelout<=1'b1;
8808: pixelout<=1'b1;
8809: pixelout<=1'b1;
8810: pixelout<=1'b1;
8811: pixelout<=1'b1;
8812: pixelout<=1'b1;
8813: pixelout<=1'b1;
8814: pixelout<=1'b1;
8815: pixelout<=1'b1;
8816: pixelout<=1'b1;
8817: pixelout<=1'b1;
8818: pixelout<=1'b1;
8819: pixelout<=1'b1;
8820: pixelout<=1'b1;
8821: pixelout<=1'b1;
8822: pixelout<=1'b0;
8823: pixelout<=1'b1;
8824: pixelout<=1'b1;
8825: pixelout<=1'b1;
8826: pixelout<=1'b1;
8827: pixelout<=1'b1;
8828: pixelout<=1'b1;
8829: pixelout<=1'b1;
8830: pixelout<=1'b1;
8831: pixelout<=1'b1;
8832: pixelout<=1'b1;
8833: pixelout<=1'b1;
8834: pixelout<=1'b1;
8835: pixelout<=1'b1;
8836: pixelout<=1'b1;
8837: pixelout<=1'b1;
8838: pixelout<=1'b1;
8839: pixelout<=1'b1;
8840: pixelout<=1'b1;
8841: pixelout<=1'b1;
8842: pixelout<=1'b1;
8843: pixelout<=1'b1;
8844: pixelout<=1'b1;
8845: pixelout<=1'b1;
8846: pixelout<=1'b1;
8847: pixelout<=1'b1;
8848: pixelout<=1'b1;
8849: pixelout<=1'b1;
8850: pixelout<=1'b1;
8851: pixelout<=1'b1;
8852: pixelout<=1'b1;
8853: pixelout<=1'b1;
8854: pixelout<=1'b1;
8855: pixelout<=1'b1;
8856: pixelout<=1'b1;
8857: pixelout<=1'b1;
8858: pixelout<=1'b1;
8859: pixelout<=1'b1;
8860: pixelout<=1'b1;
8861: pixelout<=1'b1;
8862: pixelout<=1'b1;
8863: pixelout<=1'b1;
8864: pixelout<=1'b1;
8865: pixelout<=1'b1;
8866: pixelout<=1'b1;
8867: pixelout<=1'b1;
8868: pixelout<=1'b1;
8869: pixelout<=1'b1;
8870: pixelout<=1'b1;
8871: pixelout<=1'b1;
8872: pixelout<=1'b1;
8873: pixelout<=1'b1;
8874: pixelout<=1'b1;
8875: pixelout<=1'b1;
8876: pixelout<=1'b1;
8877: pixelout<=1'b1;
8878: pixelout<=1'b1;
8879: pixelout<=1'b1;
8880: pixelout<=1'b1;
8881: pixelout<=1'b1;
8882: pixelout<=1'b1;
8883: pixelout<=1'b1;
8884: pixelout<=1'b1;
8885: pixelout<=1'b1;
8886: pixelout<=1'b1;
8887: pixelout<=1'b1;
8888: pixelout<=1'b1;
8889: pixelout<=1'b1;
8890: pixelout<=1'b1;
8891: pixelout<=1'b1;
8892: pixelout<=1'b1;
8893: pixelout<=1'b1;
8894: pixelout<=1'b1;
8895: pixelout<=1'b1;
8896: pixelout<=1'b1;
8897: pixelout<=1'b1;
8898: pixelout<=1'b1;
8899: pixelout<=1'b1;
8900: pixelout<=1'b1;
8901: pixelout<=1'b1;
8902: pixelout<=1'b1;
8903: pixelout<=1'b1;
8904: pixelout<=1'b1;
8905: pixelout<=1'b1;
8906: pixelout<=1'b1;
8907: pixelout<=1'b1;
8908: pixelout<=1'b1;
8909: pixelout<=1'b1;
8910: pixelout<=1'b1;
8911: pixelout<=1'b1;
8912: pixelout<=1'b1;
8913: pixelout<=1'b1;
8914: pixelout<=1'b1;
8915: pixelout<=1'b1;
8916: pixelout<=1'b1;
8917: pixelout<=1'b1;
8918: pixelout<=1'b1;
8919: pixelout<=1'b1;
8920: pixelout<=1'b1;
8921: pixelout<=1'b1;
8922: pixelout<=1'b1;
8923: pixelout<=1'b1;
8924: pixelout<=1'b1;
8925: pixelout<=1'b1;
8926: pixelout<=1'b1;
8927: pixelout<=1'b1;
8928: pixelout<=1'b1;
8929: pixelout<=1'b1;
8930: pixelout<=1'b1;
8931: pixelout<=1'b1;
8932: pixelout<=1'b1;
8933: pixelout<=1'b1;
8934: pixelout<=1'b1;
8935: pixelout<=1'b1;
8936: pixelout<=1'b0;
8937: pixelout<=1'b1;
8938: pixelout<=1'b1;
8939: pixelout<=1'b1;
8940: pixelout<=1'b0;
8941: pixelout<=1'b1;
8942: pixelout<=1'b0;
8943: pixelout<=1'b1;
8944: pixelout<=1'b1;
8945: pixelout<=1'b0;
8946: pixelout<=1'b1;
8947: pixelout<=1'b1;
8948: pixelout<=1'b1;
8949: pixelout<=1'b1;
8950: pixelout<=1'b1;
8951: pixelout<=1'b1;
8952: pixelout<=1'b0;
8953: pixelout<=1'b1;
8954: pixelout<=1'b1;
8955: pixelout<=1'b1;
8956: pixelout<=1'b0;
8957: pixelout<=1'b1;
8958: pixelout<=1'b1;
8959: pixelout<=1'b1;
8960: pixelout<=1'b0;
8961: pixelout<=1'b1;
8962: pixelout<=1'b0;
8963: pixelout<=1'b1;
8964: pixelout<=1'b1;
8965: pixelout<=1'b1;
8966: pixelout<=1'b0;
8967: pixelout<=1'b1;
8968: pixelout<=1'b0;
8969: pixelout<=1'b1;
8970: pixelout<=1'b1;
8971: pixelout<=1'b0;
8972: pixelout<=1'b1;
8973: pixelout<=1'b1;
8974: pixelout<=1'b1;
8975: pixelout<=1'b0;
8976: pixelout<=1'b1;
8977: pixelout<=1'b1;
8978: pixelout<=1'b1;
8979: pixelout<=1'b1;
8980: pixelout<=1'b1;
8981: pixelout<=1'b1;
8982: pixelout<=1'b0;
8983: pixelout<=1'b1;
8984: pixelout<=1'b1;
8985: pixelout<=1'b1;
8986: pixelout<=1'b1;
8987: pixelout<=1'b1;
8988: pixelout<=1'b0;
8989: pixelout<=1'b1;
8990: pixelout<=1'b0;
8991: pixelout<=1'b1;
8992: pixelout<=1'b1;
8993: pixelout<=1'b0;
8994: pixelout<=1'b1;
8995: pixelout<=1'b0;
8996: pixelout<=1'b1;
8997: pixelout<=1'b1;
8998: pixelout<=1'b1;
8999: pixelout<=1'b1;
9000: pixelout<=1'b1;
9001: pixelout<=1'b1;
9002: pixelout<=1'b1;
9003: pixelout<=1'b1;
9004: pixelout<=1'b1;
9005: pixelout<=1'b1;
9006: pixelout<=1'b1;
9007: pixelout<=1'b0;
9008: pixelout<=1'b0;
9009: pixelout<=1'b0;
9010: pixelout<=1'b0;
9011: pixelout<=1'b1;
9012: pixelout<=1'b1;
9013: pixelout<=1'b0;
9014: pixelout<=1'b0;
9015: pixelout<=1'b1;
9016: pixelout<=1'b1;
9017: pixelout<=1'b1;
9018: pixelout<=1'b0;
9019: pixelout<=1'b1;
9020: pixelout<=1'b1;
9021: pixelout<=1'b1;
9022: pixelout<=1'b1;
9023: pixelout<=1'b1;
9024: pixelout<=1'b1;
9025: pixelout<=1'b1;
9026: pixelout<=1'b1;
9027: pixelout<=1'b1;
9028: pixelout<=1'b0;
9029: pixelout<=1'b1;
9030: pixelout<=1'b0;
9031: pixelout<=1'b1;
9032: pixelout<=1'b1;
9033: pixelout<=1'b1;
9034: pixelout<=1'b0;
9035: pixelout<=1'b1;
9036: pixelout<=1'b0;
9037: pixelout<=1'b1;
9038: pixelout<=1'b1;
9039: pixelout<=1'b1;
9040: pixelout<=1'b0;
9041: pixelout<=1'b1;
9042: pixelout<=1'b1;
9043: pixelout<=1'b0;
9044: pixelout<=1'b1;
9045: pixelout<=1'b1;
9046: pixelout<=1'b1;
9047: pixelout<=1'b1;
9048: pixelout<=1'b1;
9049: pixelout<=1'b1;
9050: pixelout<=1'b1;
9051: pixelout<=1'b1;
9052: pixelout<=1'b1;
9053: pixelout<=1'b1;
9054: pixelout<=1'b1;
9055: pixelout<=1'b1;
9056: pixelout<=1'b1;
9057: pixelout<=1'b1;
9058: pixelout<=1'b1;
9059: pixelout<=1'b1;
9060: pixelout<=1'b1;
9061: pixelout<=1'b1;
9062: pixelout<=1'b0;
9063: pixelout<=1'b1;
9064: pixelout<=1'b1;
9065: pixelout<=1'b1;
9066: pixelout<=1'b1;
9067: pixelout<=1'b1;
9068: pixelout<=1'b1;
9069: pixelout<=1'b1;
9070: pixelout<=1'b1;
9071: pixelout<=1'b1;
9072: pixelout<=1'b1;
9073: pixelout<=1'b1;
9074: pixelout<=1'b1;
9075: pixelout<=1'b1;
9076: pixelout<=1'b1;
9077: pixelout<=1'b1;
9078: pixelout<=1'b1;
9079: pixelout<=1'b1;
9080: pixelout<=1'b1;
9081: pixelout<=1'b1;
9082: pixelout<=1'b1;
9083: pixelout<=1'b1;
9084: pixelout<=1'b1;
9085: pixelout<=1'b1;
9086: pixelout<=1'b1;
9087: pixelout<=1'b1;
9088: pixelout<=1'b1;
9089: pixelout<=1'b1;
9090: pixelout<=1'b1;
9091: pixelout<=1'b1;
9092: pixelout<=1'b1;
9093: pixelout<=1'b1;
9094: pixelout<=1'b1;
9095: pixelout<=1'b1;
9096: pixelout<=1'b1;
9097: pixelout<=1'b1;
9098: pixelout<=1'b1;
9099: pixelout<=1'b1;
9100: pixelout<=1'b1;
9101: pixelout<=1'b1;
9102: pixelout<=1'b1;
9103: pixelout<=1'b1;
9104: pixelout<=1'b1;
9105: pixelout<=1'b1;
9106: pixelout<=1'b1;
9107: pixelout<=1'b1;
9108: pixelout<=1'b1;
9109: pixelout<=1'b1;
9110: pixelout<=1'b1;
9111: pixelout<=1'b1;
9112: pixelout<=1'b1;
9113: pixelout<=1'b1;
9114: pixelout<=1'b1;
9115: pixelout<=1'b1;
9116: pixelout<=1'b1;
9117: pixelout<=1'b1;
9118: pixelout<=1'b1;
9119: pixelout<=1'b1;
9120: pixelout<=1'b1;
9121: pixelout<=1'b1;
9122: pixelout<=1'b1;
9123: pixelout<=1'b1;
9124: pixelout<=1'b1;
9125: pixelout<=1'b1;
9126: pixelout<=1'b1;
9127: pixelout<=1'b1;
9128: pixelout<=1'b1;
9129: pixelout<=1'b1;
9130: pixelout<=1'b1;
9131: pixelout<=1'b1;
9132: pixelout<=1'b1;
9133: pixelout<=1'b1;
9134: pixelout<=1'b1;
9135: pixelout<=1'b1;
9136: pixelout<=1'b1;
9137: pixelout<=1'b1;
9138: pixelout<=1'b1;
9139: pixelout<=1'b1;
9140: pixelout<=1'b1;
9141: pixelout<=1'b1;
9142: pixelout<=1'b1;
9143: pixelout<=1'b1;
9144: pixelout<=1'b1;
9145: pixelout<=1'b1;
9146: pixelout<=1'b1;
9147: pixelout<=1'b1;
9148: pixelout<=1'b1;
9149: pixelout<=1'b1;
9150: pixelout<=1'b1;
9151: pixelout<=1'b1;
9152: pixelout<=1'b1;
9153: pixelout<=1'b1;
9154: pixelout<=1'b1;
9155: pixelout<=1'b1;
9156: pixelout<=1'b1;
9157: pixelout<=1'b1;
9158: pixelout<=1'b1;
9159: pixelout<=1'b1;
9160: pixelout<=1'b1;
9161: pixelout<=1'b1;
9162: pixelout<=1'b1;
9163: pixelout<=1'b1;
9164: pixelout<=1'b1;
9165: pixelout<=1'b1;
9166: pixelout<=1'b1;
9167: pixelout<=1'b1;
9168: pixelout<=1'b1;
9169: pixelout<=1'b1;
9170: pixelout<=1'b1;
9171: pixelout<=1'b1;
9172: pixelout<=1'b1;
9173: pixelout<=1'b1;
9174: pixelout<=1'b1;
9175: pixelout<=1'b1;
9176: pixelout<=1'b0;
9177: pixelout<=1'b1;
9178: pixelout<=1'b1;
9179: pixelout<=1'b1;
9180: pixelout<=1'b0;
9181: pixelout<=1'b1;
9182: pixelout<=1'b0;
9183: pixelout<=1'b1;
9184: pixelout<=1'b1;
9185: pixelout<=1'b0;
9186: pixelout<=1'b1;
9187: pixelout<=1'b1;
9188: pixelout<=1'b1;
9189: pixelout<=1'b1;
9190: pixelout<=1'b1;
9191: pixelout<=1'b1;
9192: pixelout<=1'b0;
9193: pixelout<=1'b1;
9194: pixelout<=1'b1;
9195: pixelout<=1'b1;
9196: pixelout<=1'b0;
9197: pixelout<=1'b1;
9198: pixelout<=1'b1;
9199: pixelout<=1'b1;
9200: pixelout<=1'b0;
9201: pixelout<=1'b1;
9202: pixelout<=1'b0;
9203: pixelout<=1'b1;
9204: pixelout<=1'b1;
9205: pixelout<=1'b1;
9206: pixelout<=1'b0;
9207: pixelout<=1'b1;
9208: pixelout<=1'b0;
9209: pixelout<=1'b1;
9210: pixelout<=1'b1;
9211: pixelout<=1'b0;
9212: pixelout<=1'b1;
9213: pixelout<=1'b1;
9214: pixelout<=1'b1;
9215: pixelout<=1'b1;
9216: pixelout<=1'b1;
9217: pixelout<=1'b1;
9218: pixelout<=1'b1;
9219: pixelout<=1'b1;
9220: pixelout<=1'b1;
9221: pixelout<=1'b1;
9222: pixelout<=1'b0;
9223: pixelout<=1'b1;
9224: pixelout<=1'b1;
9225: pixelout<=1'b1;
9226: pixelout<=1'b1;
9227: pixelout<=1'b1;
9228: pixelout<=1'b0;
9229: pixelout<=1'b1;
9230: pixelout<=1'b0;
9231: pixelout<=1'b1;
9232: pixelout<=1'b1;
9233: pixelout<=1'b0;
9234: pixelout<=1'b1;
9235: pixelout<=1'b0;
9236: pixelout<=1'b1;
9237: pixelout<=1'b1;
9238: pixelout<=1'b1;
9239: pixelout<=1'b1;
9240: pixelout<=1'b1;
9241: pixelout<=1'b1;
9242: pixelout<=1'b1;
9243: pixelout<=1'b1;
9244: pixelout<=1'b1;
9245: pixelout<=1'b1;
9246: pixelout<=1'b1;
9247: pixelout<=1'b0;
9248: pixelout<=1'b1;
9249: pixelout<=1'b1;
9250: pixelout<=1'b1;
9251: pixelout<=1'b1;
9252: pixelout<=1'b1;
9253: pixelout<=1'b0;
9254: pixelout<=1'b1;
9255: pixelout<=1'b1;
9256: pixelout<=1'b1;
9257: pixelout<=1'b1;
9258: pixelout<=1'b0;
9259: pixelout<=1'b1;
9260: pixelout<=1'b1;
9261: pixelout<=1'b1;
9262: pixelout<=1'b1;
9263: pixelout<=1'b1;
9264: pixelout<=1'b1;
9265: pixelout<=1'b1;
9266: pixelout<=1'b1;
9267: pixelout<=1'b1;
9268: pixelout<=1'b0;
9269: pixelout<=1'b1;
9270: pixelout<=1'b0;
9271: pixelout<=1'b0;
9272: pixelout<=1'b0;
9273: pixelout<=1'b0;
9274: pixelout<=1'b0;
9275: pixelout<=1'b1;
9276: pixelout<=1'b0;
9277: pixelout<=1'b1;
9278: pixelout<=1'b1;
9279: pixelout<=1'b1;
9280: pixelout<=1'b1;
9281: pixelout<=1'b1;
9282: pixelout<=1'b1;
9283: pixelout<=1'b0;
9284: pixelout<=1'b1;
9285: pixelout<=1'b1;
9286: pixelout<=1'b1;
9287: pixelout<=1'b1;
9288: pixelout<=1'b1;
9289: pixelout<=1'b1;
9290: pixelout<=1'b1;
9291: pixelout<=1'b1;
9292: pixelout<=1'b1;
9293: pixelout<=1'b1;
9294: pixelout<=1'b1;
9295: pixelout<=1'b1;
9296: pixelout<=1'b1;
9297: pixelout<=1'b1;
9298: pixelout<=1'b0;
9299: pixelout<=1'b0;
9300: pixelout<=1'b1;
9301: pixelout<=1'b1;
9302: pixelout<=1'b0;
9303: pixelout<=1'b1;
9304: pixelout<=1'b1;
9305: pixelout<=1'b1;
9306: pixelout<=1'b1;
9307: pixelout<=1'b1;
9308: pixelout<=1'b1;
9309: pixelout<=1'b1;
9310: pixelout<=1'b1;
9311: pixelout<=1'b1;
9312: pixelout<=1'b1;
9313: pixelout<=1'b1;
9314: pixelout<=1'b1;
9315: pixelout<=1'b1;
9316: pixelout<=1'b1;
9317: pixelout<=1'b1;
9318: pixelout<=1'b1;
9319: pixelout<=1'b1;
9320: pixelout<=1'b1;
9321: pixelout<=1'b1;
9322: pixelout<=1'b1;
9323: pixelout<=1'b1;
9324: pixelout<=1'b1;
9325: pixelout<=1'b1;
9326: pixelout<=1'b1;
9327: pixelout<=1'b1;
9328: pixelout<=1'b1;
9329: pixelout<=1'b1;
9330: pixelout<=1'b1;
9331: pixelout<=1'b1;
9332: pixelout<=1'b1;
9333: pixelout<=1'b1;
9334: pixelout<=1'b1;
9335: pixelout<=1'b1;
9336: pixelout<=1'b1;
9337: pixelout<=1'b1;
9338: pixelout<=1'b1;
9339: pixelout<=1'b1;
9340: pixelout<=1'b1;
9341: pixelout<=1'b1;
9342: pixelout<=1'b1;
9343: pixelout<=1'b1;
9344: pixelout<=1'b1;
9345: pixelout<=1'b1;
9346: pixelout<=1'b1;
9347: pixelout<=1'b1;
9348: pixelout<=1'b1;
9349: pixelout<=1'b1;
9350: pixelout<=1'b1;
9351: pixelout<=1'b1;
9352: pixelout<=1'b1;
9353: pixelout<=1'b1;
9354: pixelout<=1'b1;
9355: pixelout<=1'b1;
9356: pixelout<=1'b1;
9357: pixelout<=1'b1;
9358: pixelout<=1'b1;
9359: pixelout<=1'b1;
9360: pixelout<=1'b1;
9361: pixelout<=1'b1;
9362: pixelout<=1'b1;
9363: pixelout<=1'b1;
9364: pixelout<=1'b1;
9365: pixelout<=1'b1;
9366: pixelout<=1'b1;
9367: pixelout<=1'b1;
9368: pixelout<=1'b1;
9369: pixelout<=1'b1;
9370: pixelout<=1'b1;
9371: pixelout<=1'b1;
9372: pixelout<=1'b1;
9373: pixelout<=1'b1;
9374: pixelout<=1'b1;
9375: pixelout<=1'b1;
9376: pixelout<=1'b1;
9377: pixelout<=1'b1;
9378: pixelout<=1'b1;
9379: pixelout<=1'b1;
9380: pixelout<=1'b1;
9381: pixelout<=1'b1;
9382: pixelout<=1'b1;
9383: pixelout<=1'b1;
9384: pixelout<=1'b1;
9385: pixelout<=1'b1;
9386: pixelout<=1'b1;
9387: pixelout<=1'b1;
9388: pixelout<=1'b1;
9389: pixelout<=1'b1;
9390: pixelout<=1'b1;
9391: pixelout<=1'b1;
9392: pixelout<=1'b1;
9393: pixelout<=1'b1;
9394: pixelout<=1'b1;
9395: pixelout<=1'b1;
9396: pixelout<=1'b1;
9397: pixelout<=1'b1;
9398: pixelout<=1'b1;
9399: pixelout<=1'b1;
9400: pixelout<=1'b1;
9401: pixelout<=1'b1;
9402: pixelout<=1'b1;
9403: pixelout<=1'b1;
9404: pixelout<=1'b1;
9405: pixelout<=1'b1;
9406: pixelout<=1'b1;
9407: pixelout<=1'b1;
9408: pixelout<=1'b1;
9409: pixelout<=1'b1;
9410: pixelout<=1'b1;
9411: pixelout<=1'b1;
9412: pixelout<=1'b1;
9413: pixelout<=1'b1;
9414: pixelout<=1'b1;
9415: pixelout<=1'b1;
9416: pixelout<=1'b0;
9417: pixelout<=1'b1;
9418: pixelout<=1'b1;
9419: pixelout<=1'b0;
9420: pixelout<=1'b0;
9421: pixelout<=1'b1;
9422: pixelout<=1'b0;
9423: pixelout<=1'b1;
9424: pixelout<=1'b1;
9425: pixelout<=1'b0;
9426: pixelout<=1'b1;
9427: pixelout<=1'b1;
9428: pixelout<=1'b1;
9429: pixelout<=1'b1;
9430: pixelout<=1'b1;
9431: pixelout<=1'b1;
9432: pixelout<=1'b0;
9433: pixelout<=1'b1;
9434: pixelout<=1'b1;
9435: pixelout<=1'b1;
9436: pixelout<=1'b0;
9437: pixelout<=1'b1;
9438: pixelout<=1'b1;
9439: pixelout<=1'b1;
9440: pixelout<=1'b0;
9441: pixelout<=1'b1;
9442: pixelout<=1'b0;
9443: pixelout<=1'b1;
9444: pixelout<=1'b1;
9445: pixelout<=1'b1;
9446: pixelout<=1'b0;
9447: pixelout<=1'b1;
9448: pixelout<=1'b0;
9449: pixelout<=1'b1;
9450: pixelout<=1'b1;
9451: pixelout<=1'b0;
9452: pixelout<=1'b1;
9453: pixelout<=1'b1;
9454: pixelout<=1'b1;
9455: pixelout<=1'b1;
9456: pixelout<=1'b1;
9457: pixelout<=1'b1;
9458: pixelout<=1'b1;
9459: pixelout<=1'b1;
9460: pixelout<=1'b1;
9461: pixelout<=1'b1;
9462: pixelout<=1'b0;
9463: pixelout<=1'b1;
9464: pixelout<=1'b1;
9465: pixelout<=1'b1;
9466: pixelout<=1'b1;
9467: pixelout<=1'b1;
9468: pixelout<=1'b0;
9469: pixelout<=1'b1;
9470: pixelout<=1'b0;
9471: pixelout<=1'b1;
9472: pixelout<=1'b1;
9473: pixelout<=1'b0;
9474: pixelout<=1'b1;
9475: pixelout<=1'b0;
9476: pixelout<=1'b1;
9477: pixelout<=1'b1;
9478: pixelout<=1'b0;
9479: pixelout<=1'b0;
9480: pixelout<=1'b1;
9481: pixelout<=1'b1;
9482: pixelout<=1'b1;
9483: pixelout<=1'b1;
9484: pixelout<=1'b1;
9485: pixelout<=1'b1;
9486: pixelout<=1'b1;
9487: pixelout<=1'b0;
9488: pixelout<=1'b1;
9489: pixelout<=1'b1;
9490: pixelout<=1'b1;
9491: pixelout<=1'b1;
9492: pixelout<=1'b1;
9493: pixelout<=1'b0;
9494: pixelout<=1'b1;
9495: pixelout<=1'b1;
9496: pixelout<=1'b1;
9497: pixelout<=1'b1;
9498: pixelout<=1'b0;
9499: pixelout<=1'b1;
9500: pixelout<=1'b1;
9501: pixelout<=1'b1;
9502: pixelout<=1'b1;
9503: pixelout<=1'b1;
9504: pixelout<=1'b1;
9505: pixelout<=1'b1;
9506: pixelout<=1'b1;
9507: pixelout<=1'b1;
9508: pixelout<=1'b0;
9509: pixelout<=1'b1;
9510: pixelout<=1'b0;
9511: pixelout<=1'b1;
9512: pixelout<=1'b1;
9513: pixelout<=1'b1;
9514: pixelout<=1'b1;
9515: pixelout<=1'b1;
9516: pixelout<=1'b0;
9517: pixelout<=1'b1;
9518: pixelout<=1'b1;
9519: pixelout<=1'b1;
9520: pixelout<=1'b0;
9521: pixelout<=1'b1;
9522: pixelout<=1'b1;
9523: pixelout<=1'b0;
9524: pixelout<=1'b1;
9525: pixelout<=1'b1;
9526: pixelout<=1'b1;
9527: pixelout<=1'b1;
9528: pixelout<=1'b1;
9529: pixelout<=1'b1;
9530: pixelout<=1'b1;
9531: pixelout<=1'b1;
9532: pixelout<=1'b1;
9533: pixelout<=1'b1;
9534: pixelout<=1'b1;
9535: pixelout<=1'b1;
9536: pixelout<=1'b1;
9537: pixelout<=1'b1;
9538: pixelout<=1'b0;
9539: pixelout<=1'b0;
9540: pixelout<=1'b1;
9541: pixelout<=1'b1;
9542: pixelout<=1'b0;
9543: pixelout<=1'b1;
9544: pixelout<=1'b1;
9545: pixelout<=1'b1;
9546: pixelout<=1'b1;
9547: pixelout<=1'b1;
9548: pixelout<=1'b1;
9549: pixelout<=1'b1;
9550: pixelout<=1'b1;
9551: pixelout<=1'b1;
9552: pixelout<=1'b1;
9553: pixelout<=1'b1;
9554: pixelout<=1'b1;
9555: pixelout<=1'b1;
9556: pixelout<=1'b1;
9557: pixelout<=1'b1;
9558: pixelout<=1'b1;
9559: pixelout<=1'b1;
9560: pixelout<=1'b1;
9561: pixelout<=1'b1;
9562: pixelout<=1'b1;
9563: pixelout<=1'b1;
9564: pixelout<=1'b1;
9565: pixelout<=1'b1;
9566: pixelout<=1'b1;
9567: pixelout<=1'b1;
9568: pixelout<=1'b1;
9569: pixelout<=1'b1;
9570: pixelout<=1'b1;
9571: pixelout<=1'b1;
9572: pixelout<=1'b1;
9573: pixelout<=1'b1;
9574: pixelout<=1'b1;
9575: pixelout<=1'b1;
9576: pixelout<=1'b1;
9577: pixelout<=1'b1;
9578: pixelout<=1'b1;
9579: pixelout<=1'b1;
9580: pixelout<=1'b1;
9581: pixelout<=1'b1;
9582: pixelout<=1'b1;
9583: pixelout<=1'b1;
9584: pixelout<=1'b1;
9585: pixelout<=1'b1;
9586: pixelout<=1'b1;
9587: pixelout<=1'b1;
9588: pixelout<=1'b1;
9589: pixelout<=1'b1;
9590: pixelout<=1'b1;
9591: pixelout<=1'b1;
9592: pixelout<=1'b1;
9593: pixelout<=1'b1;
9594: pixelout<=1'b1;
9595: pixelout<=1'b1;
9596: pixelout<=1'b1;
9597: pixelout<=1'b1;
9598: pixelout<=1'b1;
9599: pixelout<=1'b1;
9600: pixelout<=1'b1;
9601: pixelout<=1'b1;
9602: pixelout<=1'b1;
9603: pixelout<=1'b1;
9604: pixelout<=1'b1;
9605: pixelout<=1'b1;
9606: pixelout<=1'b1;
9607: pixelout<=1'b1;
9608: pixelout<=1'b1;
9609: pixelout<=1'b1;
9610: pixelout<=1'b1;
9611: pixelout<=1'b1;
9612: pixelout<=1'b1;
9613: pixelout<=1'b1;
9614: pixelout<=1'b1;
9615: pixelout<=1'b1;
9616: pixelout<=1'b1;
9617: pixelout<=1'b1;
9618: pixelout<=1'b1;
9619: pixelout<=1'b1;
9620: pixelout<=1'b1;
9621: pixelout<=1'b1;
9622: pixelout<=1'b1;
9623: pixelout<=1'b1;
9624: pixelout<=1'b1;
9625: pixelout<=1'b1;
9626: pixelout<=1'b1;
9627: pixelout<=1'b1;
9628: pixelout<=1'b1;
9629: pixelout<=1'b1;
9630: pixelout<=1'b1;
9631: pixelout<=1'b1;
9632: pixelout<=1'b1;
9633: pixelout<=1'b1;
9634: pixelout<=1'b1;
9635: pixelout<=1'b1;
9636: pixelout<=1'b1;
9637: pixelout<=1'b1;
9638: pixelout<=1'b1;
9639: pixelout<=1'b1;
9640: pixelout<=1'b1;
9641: pixelout<=1'b1;
9642: pixelout<=1'b1;
9643: pixelout<=1'b1;
9644: pixelout<=1'b1;
9645: pixelout<=1'b1;
9646: pixelout<=1'b1;
9647: pixelout<=1'b1;
9648: pixelout<=1'b1;
9649: pixelout<=1'b1;
9650: pixelout<=1'b1;
9651: pixelout<=1'b1;
9652: pixelout<=1'b1;
9653: pixelout<=1'b1;
9654: pixelout<=1'b1;
9655: pixelout<=1'b1;
9656: pixelout<=1'b1;
9657: pixelout<=1'b0;
9658: pixelout<=1'b0;
9659: pixelout<=1'b1;
9660: pixelout<=1'b0;
9661: pixelout<=1'b1;
9662: pixelout<=1'b0;
9663: pixelout<=1'b1;
9664: pixelout<=1'b1;
9665: pixelout<=1'b0;
9666: pixelout<=1'b1;
9667: pixelout<=1'b1;
9668: pixelout<=1'b1;
9669: pixelout<=1'b0;
9670: pixelout<=1'b0;
9671: pixelout<=1'b0;
9672: pixelout<=1'b0;
9673: pixelout<=1'b1;
9674: pixelout<=1'b1;
9675: pixelout<=1'b1;
9676: pixelout<=1'b1;
9677: pixelout<=1'b0;
9678: pixelout<=1'b0;
9679: pixelout<=1'b0;
9680: pixelout<=1'b0;
9681: pixelout<=1'b1;
9682: pixelout<=1'b1;
9683: pixelout<=1'b0;
9684: pixelout<=1'b0;
9685: pixelout<=1'b0;
9686: pixelout<=1'b1;
9687: pixelout<=1'b1;
9688: pixelout<=1'b1;
9689: pixelout<=1'b0;
9690: pixelout<=1'b0;
9691: pixelout<=1'b1;
9692: pixelout<=1'b1;
9693: pixelout<=1'b1;
9694: pixelout<=1'b1;
9695: pixelout<=1'b1;
9696: pixelout<=1'b1;
9697: pixelout<=1'b1;
9698: pixelout<=1'b1;
9699: pixelout<=1'b1;
9700: pixelout<=1'b1;
9701: pixelout<=1'b1;
9702: pixelout<=1'b0;
9703: pixelout<=1'b1;
9704: pixelout<=1'b1;
9705: pixelout<=1'b1;
9706: pixelout<=1'b1;
9707: pixelout<=1'b1;
9708: pixelout<=1'b0;
9709: pixelout<=1'b1;
9710: pixelout<=1'b0;
9711: pixelout<=1'b1;
9712: pixelout<=1'b1;
9713: pixelout<=1'b0;
9714: pixelout<=1'b1;
9715: pixelout<=1'b1;
9716: pixelout<=1'b0;
9717: pixelout<=1'b0;
9718: pixelout<=1'b1;
9719: pixelout<=1'b1;
9720: pixelout<=1'b1;
9721: pixelout<=1'b1;
9722: pixelout<=1'b1;
9723: pixelout<=1'b1;
9724: pixelout<=1'b1;
9725: pixelout<=1'b1;
9726: pixelout<=1'b1;
9727: pixelout<=1'b0;
9728: pixelout<=1'b1;
9729: pixelout<=1'b1;
9730: pixelout<=1'b1;
9731: pixelout<=1'b1;
9732: pixelout<=1'b1;
9733: pixelout<=1'b0;
9734: pixelout<=1'b1;
9735: pixelout<=1'b1;
9736: pixelout<=1'b1;
9737: pixelout<=1'b1;
9738: pixelout<=1'b1;
9739: pixelout<=1'b0;
9740: pixelout<=1'b0;
9741: pixelout<=1'b0;
9742: pixelout<=1'b1;
9743: pixelout<=1'b1;
9744: pixelout<=1'b1;
9745: pixelout<=1'b1;
9746: pixelout<=1'b1;
9747: pixelout<=1'b1;
9748: pixelout<=1'b0;
9749: pixelout<=1'b1;
9750: pixelout<=1'b1;
9751: pixelout<=1'b0;
9752: pixelout<=1'b0;
9753: pixelout<=1'b0;
9754: pixelout<=1'b0;
9755: pixelout<=1'b1;
9756: pixelout<=1'b1;
9757: pixelout<=1'b0;
9758: pixelout<=1'b0;
9759: pixelout<=1'b0;
9760: pixelout<=1'b1;
9761: pixelout<=1'b1;
9762: pixelout<=1'b1;
9763: pixelout<=1'b0;
9764: pixelout<=1'b0;
9765: pixelout<=1'b0;
9766: pixelout<=1'b1;
9767: pixelout<=1'b1;
9768: pixelout<=1'b1;
9769: pixelout<=1'b1;
9770: pixelout<=1'b1;
9771: pixelout<=1'b1;
9772: pixelout<=1'b1;
9773: pixelout<=1'b1;
9774: pixelout<=1'b1;
9775: pixelout<=1'b1;
9776: pixelout<=1'b1;
9777: pixelout<=1'b1;
9778: pixelout<=1'b1;
9779: pixelout<=1'b0;
9780: pixelout<=1'b1;
9781: pixelout<=1'b0;
9782: pixelout<=1'b1;
9783: pixelout<=1'b1;
9784: pixelout<=1'b1;
9785: pixelout<=1'b1;
9786: pixelout<=1'b1;
9787: pixelout<=1'b1;
9788: pixelout<=1'b1;
9789: pixelout<=1'b1;
9790: pixelout<=1'b1;
9791: pixelout<=1'b1;
9792: pixelout<=1'b1;
9793: pixelout<=1'b1;
9794: pixelout<=1'b1;
9795: pixelout<=1'b1;
9796: pixelout<=1'b1;
9797: pixelout<=1'b1;
9798: pixelout<=1'b1;
9799: pixelout<=1'b1;
9800: pixelout<=1'b1;
9801: pixelout<=1'b1;
9802: pixelout<=1'b1;
9803: pixelout<=1'b1;
9804: pixelout<=1'b1;
9805: pixelout<=1'b1;
9806: pixelout<=1'b1;
9807: pixelout<=1'b1;
9808: pixelout<=1'b1;
9809: pixelout<=1'b1;
9810: pixelout<=1'b1;
9811: pixelout<=1'b1;
9812: pixelout<=1'b1;
9813: pixelout<=1'b1;
9814: pixelout<=1'b1;
9815: pixelout<=1'b1;
9816: pixelout<=1'b1;
9817: pixelout<=1'b1;
9818: pixelout<=1'b1;
9819: pixelout<=1'b1;
9820: pixelout<=1'b1;
9821: pixelout<=1'b1;
9822: pixelout<=1'b1;
9823: pixelout<=1'b1;
9824: pixelout<=1'b1;
9825: pixelout<=1'b1;
9826: pixelout<=1'b1;
9827: pixelout<=1'b1;
9828: pixelout<=1'b1;
9829: pixelout<=1'b1;
9830: pixelout<=1'b1;
9831: pixelout<=1'b1;
9832: pixelout<=1'b1;
9833: pixelout<=1'b1;
9834: pixelout<=1'b1;
9835: pixelout<=1'b1;
9836: pixelout<=1'b1;
9837: pixelout<=1'b1;
9838: pixelout<=1'b1;
9839: pixelout<=1'b1;
9840: pixelout<=1'b1;
9841: pixelout<=1'b1;
9842: pixelout<=1'b1;
9843: pixelout<=1'b1;
9844: pixelout<=1'b1;
9845: pixelout<=1'b1;
9846: pixelout<=1'b1;
9847: pixelout<=1'b1;
9848: pixelout<=1'b1;
9849: pixelout<=1'b1;
9850: pixelout<=1'b1;
9851: pixelout<=1'b1;
9852: pixelout<=1'b1;
9853: pixelout<=1'b1;
9854: pixelout<=1'b1;
9855: pixelout<=1'b1;
9856: pixelout<=1'b1;
9857: pixelout<=1'b1;
9858: pixelout<=1'b1;
9859: pixelout<=1'b1;
9860: pixelout<=1'b1;
9861: pixelout<=1'b1;
9862: pixelout<=1'b1;
9863: pixelout<=1'b1;
9864: pixelout<=1'b1;
9865: pixelout<=1'b1;
9866: pixelout<=1'b1;
9867: pixelout<=1'b1;
9868: pixelout<=1'b1;
9869: pixelout<=1'b1;
9870: pixelout<=1'b1;
9871: pixelout<=1'b1;
9872: pixelout<=1'b1;
9873: pixelout<=1'b1;
9874: pixelout<=1'b1;
9875: pixelout<=1'b1;
9876: pixelout<=1'b1;
9877: pixelout<=1'b1;
9878: pixelout<=1'b1;
9879: pixelout<=1'b1;
9880: pixelout<=1'b1;
9881: pixelout<=1'b1;
9882: pixelout<=1'b1;
9883: pixelout<=1'b1;
9884: pixelout<=1'b1;
9885: pixelout<=1'b1;
9886: pixelout<=1'b1;
9887: pixelout<=1'b1;
9888: pixelout<=1'b1;
9889: pixelout<=1'b1;
9890: pixelout<=1'b1;
9891: pixelout<=1'b1;
9892: pixelout<=1'b1;
9893: pixelout<=1'b1;
9894: pixelout<=1'b1;
9895: pixelout<=1'b1;
9896: pixelout<=1'b1;
9897: pixelout<=1'b1;
9898: pixelout<=1'b1;
9899: pixelout<=1'b1;
9900: pixelout<=1'b1;
9901: pixelout<=1'b1;
9902: pixelout<=1'b1;
9903: pixelout<=1'b1;
9904: pixelout<=1'b1;
9905: pixelout<=1'b1;
9906: pixelout<=1'b1;
9907: pixelout<=1'b1;
9908: pixelout<=1'b1;
9909: pixelout<=1'b1;
9910: pixelout<=1'b1;
9911: pixelout<=1'b1;
9912: pixelout<=1'b1;
9913: pixelout<=1'b1;
9914: pixelout<=1'b1;
9915: pixelout<=1'b1;
9916: pixelout<=1'b1;
9917: pixelout<=1'b1;
9918: pixelout<=1'b1;
9919: pixelout<=1'b1;
9920: pixelout<=1'b0;
9921: pixelout<=1'b1;
9922: pixelout<=1'b1;
9923: pixelout<=1'b1;
9924: pixelout<=1'b1;
9925: pixelout<=1'b1;
9926: pixelout<=1'b1;
9927: pixelout<=1'b1;
9928: pixelout<=1'b1;
9929: pixelout<=1'b1;
9930: pixelout<=1'b1;
9931: pixelout<=1'b1;
9932: pixelout<=1'b1;
9933: pixelout<=1'b1;
9934: pixelout<=1'b1;
9935: pixelout<=1'b1;
9936: pixelout<=1'b1;
9937: pixelout<=1'b1;
9938: pixelout<=1'b1;
9939: pixelout<=1'b1;
9940: pixelout<=1'b1;
9941: pixelout<=1'b1;
9942: pixelout<=1'b1;
9943: pixelout<=1'b1;
9944: pixelout<=1'b1;
9945: pixelout<=1'b1;
9946: pixelout<=1'b1;
9947: pixelout<=1'b1;
9948: pixelout<=1'b1;
9949: pixelout<=1'b1;
9950: pixelout<=1'b1;
9951: pixelout<=1'b1;
9952: pixelout<=1'b1;
9953: pixelout<=1'b1;
9954: pixelout<=1'b1;
9955: pixelout<=1'b1;
9956: pixelout<=1'b1;
9957: pixelout<=1'b1;
9958: pixelout<=1'b1;
9959: pixelout<=1'b1;
9960: pixelout<=1'b1;
9961: pixelout<=1'b1;
9962: pixelout<=1'b1;
9963: pixelout<=1'b1;
9964: pixelout<=1'b1;
9965: pixelout<=1'b1;
9966: pixelout<=1'b1;
9967: pixelout<=1'b1;
9968: pixelout<=1'b1;
9969: pixelout<=1'b1;
9970: pixelout<=1'b1;
9971: pixelout<=1'b1;
9972: pixelout<=1'b1;
9973: pixelout<=1'b1;
9974: pixelout<=1'b1;
9975: pixelout<=1'b1;
9976: pixelout<=1'b1;
9977: pixelout<=1'b1;
9978: pixelout<=1'b1;
9979: pixelout<=1'b1;
9980: pixelout<=1'b1;
9981: pixelout<=1'b1;
9982: pixelout<=1'b1;
9983: pixelout<=1'b1;
9984: pixelout<=1'b1;
9985: pixelout<=1'b1;
9986: pixelout<=1'b1;
9987: pixelout<=1'b1;
9988: pixelout<=1'b0;
9989: pixelout<=1'b1;
9990: pixelout<=1'b1;
9991: pixelout<=1'b1;
9992: pixelout<=1'b1;
9993: pixelout<=1'b1;
9994: pixelout<=1'b1;
9995: pixelout<=1'b1;
9996: pixelout<=1'b1;
9997: pixelout<=1'b1;
9998: pixelout<=1'b1;
9999: pixelout<=1'b1;
10000: pixelout<=1'b1;
10001: pixelout<=1'b1;
10002: pixelout<=1'b1;
10003: pixelout<=1'b1;
10004: pixelout<=1'b1;
10005: pixelout<=1'b1;
10006: pixelout<=1'b1;
10007: pixelout<=1'b1;
10008: pixelout<=1'b1;
10009: pixelout<=1'b1;
10010: pixelout<=1'b1;
10011: pixelout<=1'b1;
10012: pixelout<=1'b1;
10013: pixelout<=1'b1;
10014: pixelout<=1'b1;
10015: pixelout<=1'b1;
10016: pixelout<=1'b1;
10017: pixelout<=1'b1;
10018: pixelout<=1'b0;
10019: pixelout<=1'b1;
10020: pixelout<=1'b1;
10021: pixelout<=1'b1;
10022: pixelout<=1'b1;
10023: pixelout<=1'b1;
10024: pixelout<=1'b1;
10025: pixelout<=1'b1;
10026: pixelout<=1'b1;
10027: pixelout<=1'b1;
10028: pixelout<=1'b1;
10029: pixelout<=1'b1;
10030: pixelout<=1'b1;
10031: pixelout<=1'b1;
10032: pixelout<=1'b1;
10033: pixelout<=1'b1;
10034: pixelout<=1'b1;
10035: pixelout<=1'b1;
10036: pixelout<=1'b1;
10037: pixelout<=1'b1;
10038: pixelout<=1'b1;
10039: pixelout<=1'b1;
10040: pixelout<=1'b1;
10041: pixelout<=1'b1;
10042: pixelout<=1'b1;
10043: pixelout<=1'b1;
10044: pixelout<=1'b1;
10045: pixelout<=1'b1;
10046: pixelout<=1'b1;
10047: pixelout<=1'b1;
10048: pixelout<=1'b1;
10049: pixelout<=1'b1;
10050: pixelout<=1'b1;
10051: pixelout<=1'b1;
10052: pixelout<=1'b1;
10053: pixelout<=1'b1;
10054: pixelout<=1'b1;
10055: pixelout<=1'b1;
10056: pixelout<=1'b1;
10057: pixelout<=1'b1;
10058: pixelout<=1'b1;
10059: pixelout<=1'b1;
10060: pixelout<=1'b1;
10061: pixelout<=1'b1;
10062: pixelout<=1'b1;
10063: pixelout<=1'b1;
10064: pixelout<=1'b1;
10065: pixelout<=1'b1;
10066: pixelout<=1'b1;
10067: pixelout<=1'b1;
10068: pixelout<=1'b1;
10069: pixelout<=1'b1;
10070: pixelout<=1'b1;
10071: pixelout<=1'b1;
10072: pixelout<=1'b1;
10073: pixelout<=1'b1;
10074: pixelout<=1'b1;
10075: pixelout<=1'b1;
10076: pixelout<=1'b1;
10077: pixelout<=1'b1;
10078: pixelout<=1'b1;
10079: pixelout<=1'b1;
10080: pixelout<=1'b1;
10081: pixelout<=1'b1;
10082: pixelout<=1'b1;
10083: pixelout<=1'b1;
10084: pixelout<=1'b1;
10085: pixelout<=1'b1;
10086: pixelout<=1'b1;
10087: pixelout<=1'b1;
10088: pixelout<=1'b1;
10089: pixelout<=1'b1;
10090: pixelout<=1'b1;
10091: pixelout<=1'b1;
10092: pixelout<=1'b1;
10093: pixelout<=1'b1;
10094: pixelout<=1'b1;
10095: pixelout<=1'b1;
10096: pixelout<=1'b1;
10097: pixelout<=1'b1;
10098: pixelout<=1'b1;
10099: pixelout<=1'b1;
10100: pixelout<=1'b1;
10101: pixelout<=1'b1;
10102: pixelout<=1'b1;
10103: pixelout<=1'b1;
10104: pixelout<=1'b1;
10105: pixelout<=1'b1;
10106: pixelout<=1'b1;
10107: pixelout<=1'b1;
10108: pixelout<=1'b1;
10109: pixelout<=1'b1;
10110: pixelout<=1'b1;
10111: pixelout<=1'b1;
10112: pixelout<=1'b1;
10113: pixelout<=1'b1;
10114: pixelout<=1'b1;
10115: pixelout<=1'b1;
10116: pixelout<=1'b1;
10117: pixelout<=1'b1;
10118: pixelout<=1'b1;
10119: pixelout<=1'b1;
10120: pixelout<=1'b1;
10121: pixelout<=1'b1;
10122: pixelout<=1'b1;
10123: pixelout<=1'b1;
10124: pixelout<=1'b1;
10125: pixelout<=1'b1;
10126: pixelout<=1'b1;
10127: pixelout<=1'b1;
10128: pixelout<=1'b1;
10129: pixelout<=1'b1;
10130: pixelout<=1'b1;
10131: pixelout<=1'b1;
10132: pixelout<=1'b1;
10133: pixelout<=1'b1;
10134: pixelout<=1'b1;
10135: pixelout<=1'b1;
10136: pixelout<=1'b1;
10137: pixelout<=1'b1;
10138: pixelout<=1'b1;
10139: pixelout<=1'b1;
10140: pixelout<=1'b1;
10141: pixelout<=1'b1;
10142: pixelout<=1'b1;
10143: pixelout<=1'b1;
10144: pixelout<=1'b1;
10145: pixelout<=1'b1;
10146: pixelout<=1'b1;
10147: pixelout<=1'b1;
10148: pixelout<=1'b1;
10149: pixelout<=1'b1;
10150: pixelout<=1'b1;
10151: pixelout<=1'b1;
10152: pixelout<=1'b1;
10153: pixelout<=1'b1;
10154: pixelout<=1'b1;
10155: pixelout<=1'b1;
10156: pixelout<=1'b0;
10157: pixelout<=1'b0;
10158: pixelout<=1'b0;
10159: pixelout<=1'b0;
10160: pixelout<=1'b1;
10161: pixelout<=1'b1;
10162: pixelout<=1'b1;
10163: pixelout<=1'b1;
10164: pixelout<=1'b1;
10165: pixelout<=1'b1;
10166: pixelout<=1'b1;
10167: pixelout<=1'b1;
10168: pixelout<=1'b1;
10169: pixelout<=1'b1;
10170: pixelout<=1'b1;
10171: pixelout<=1'b1;
10172: pixelout<=1'b1;
10173: pixelout<=1'b1;
10174: pixelout<=1'b1;
10175: pixelout<=1'b1;
10176: pixelout<=1'b1;
10177: pixelout<=1'b1;
10178: pixelout<=1'b1;
10179: pixelout<=1'b1;
10180: pixelout<=1'b1;
10181: pixelout<=1'b1;
10182: pixelout<=1'b1;
10183: pixelout<=1'b1;
10184: pixelout<=1'b1;
10185: pixelout<=1'b1;
10186: pixelout<=1'b1;
10187: pixelout<=1'b1;
10188: pixelout<=1'b1;
10189: pixelout<=1'b1;
10190: pixelout<=1'b1;
10191: pixelout<=1'b1;
10192: pixelout<=1'b1;
10193: pixelout<=1'b1;
10194: pixelout<=1'b1;
10195: pixelout<=1'b1;
10196: pixelout<=1'b1;
10197: pixelout<=1'b1;
10198: pixelout<=1'b1;
10199: pixelout<=1'b1;
10200: pixelout<=1'b1;
10201: pixelout<=1'b1;
10202: pixelout<=1'b1;
10203: pixelout<=1'b1;
10204: pixelout<=1'b1;
10205: pixelout<=1'b1;
10206: pixelout<=1'b1;
10207: pixelout<=1'b1;
10208: pixelout<=1'b1;
10209: pixelout<=1'b1;
10210: pixelout<=1'b1;
10211: pixelout<=1'b1;
10212: pixelout<=1'b1;
10213: pixelout<=1'b1;
10214: pixelout<=1'b1;
10215: pixelout<=1'b1;
10216: pixelout<=1'b1;
10217: pixelout<=1'b1;
10218: pixelout<=1'b1;
10219: pixelout<=1'b1;
10220: pixelout<=1'b1;
10221: pixelout<=1'b1;
10222: pixelout<=1'b1;
10223: pixelout<=1'b1;
10224: pixelout<=1'b1;
10225: pixelout<=1'b1;
10226: pixelout<=1'b0;
10227: pixelout<=1'b0;
10228: pixelout<=1'b1;
10229: pixelout<=1'b1;
10230: pixelout<=1'b1;
10231: pixelout<=1'b1;
10232: pixelout<=1'b1;
10233: pixelout<=1'b1;
10234: pixelout<=1'b1;
10235: pixelout<=1'b1;
10236: pixelout<=1'b1;
10237: pixelout<=1'b1;
10238: pixelout<=1'b1;
10239: pixelout<=1'b1;
10240: pixelout<=1'b1;
10241: pixelout<=1'b1;
10242: pixelout<=1'b1;
10243: pixelout<=1'b1;
10244: pixelout<=1'b1;
10245: pixelout<=1'b1;
10246: pixelout<=1'b1;
10247: pixelout<=1'b1;
10248: pixelout<=1'b1;
10249: pixelout<=1'b1;
10250: pixelout<=1'b1;
10251: pixelout<=1'b1;
10252: pixelout<=1'b1;
10253: pixelout<=1'b1;
10254: pixelout<=1'b1;
10255: pixelout<=1'b1;
10256: pixelout<=1'b1;
10257: pixelout<=1'b1;
10258: pixelout<=1'b1;
10259: pixelout<=1'b1;
10260: pixelout<=1'b1;
10261: pixelout<=1'b1;
10262: pixelout<=1'b1;
10263: pixelout<=1'b1;
10264: pixelout<=1'b1;
10265: pixelout<=1'b1;
10266: pixelout<=1'b1;
10267: pixelout<=1'b1;
10268: pixelout<=1'b1;
10269: pixelout<=1'b1;
10270: pixelout<=1'b1;
10271: pixelout<=1'b1;
10272: pixelout<=1'b1;
10273: pixelout<=1'b1;
10274: pixelout<=1'b1;
10275: pixelout<=1'b1;
10276: pixelout<=1'b1;
10277: pixelout<=1'b1;
10278: pixelout<=1'b1;
10279: pixelout<=1'b1;
10280: pixelout<=1'b1;
10281: pixelout<=1'b1;
10282: pixelout<=1'b1;
10283: pixelout<=1'b1;
10284: pixelout<=1'b1;
10285: pixelout<=1'b1;
10286: pixelout<=1'b1;
10287: pixelout<=1'b1;
10288: pixelout<=1'b1;
10289: pixelout<=1'b1;
10290: pixelout<=1'b1;
10291: pixelout<=1'b1;
10292: pixelout<=1'b1;
10293: pixelout<=1'b1;
10294: pixelout<=1'b1;
10295: pixelout<=1'b1;
10296: pixelout<=1'b1;
10297: pixelout<=1'b1;
10298: pixelout<=1'b1;
10299: pixelout<=1'b1;
10300: pixelout<=1'b1;
10301: pixelout<=1'b1;
10302: pixelout<=1'b1;
10303: pixelout<=1'b1;
10304: pixelout<=1'b1;
10305: pixelout<=1'b1;
10306: pixelout<=1'b1;
10307: pixelout<=1'b1;
10308: pixelout<=1'b1;
10309: pixelout<=1'b1;
10310: pixelout<=1'b1;
10311: pixelout<=1'b1;
10312: pixelout<=1'b1;
10313: pixelout<=1'b1;
10314: pixelout<=1'b1;
10315: pixelout<=1'b1;
10316: pixelout<=1'b1;
10317: pixelout<=1'b1;
10318: pixelout<=1'b1;
10319: pixelout<=1'b1;
10320: pixelout<=1'b1;
10321: pixelout<=1'b1;
10322: pixelout<=1'b1;
10323: pixelout<=1'b1;
10324: pixelout<=1'b1;
10325: pixelout<=1'b1;
10326: pixelout<=1'b1;
10327: pixelout<=1'b1;
10328: pixelout<=1'b1;
10329: pixelout<=1'b1;
10330: pixelout<=1'b1;
10331: pixelout<=1'b1;
10332: pixelout<=1'b1;
10333: pixelout<=1'b1;
10334: pixelout<=1'b1;
10335: pixelout<=1'b1;
10336: pixelout<=1'b1;
10337: pixelout<=1'b1;
10338: pixelout<=1'b1;
10339: pixelout<=1'b1;
10340: pixelout<=1'b1;
10341: pixelout<=1'b1;
10342: pixelout<=1'b1;
10343: pixelout<=1'b1;
10344: pixelout<=1'b1;
10345: pixelout<=1'b1;
10346: pixelout<=1'b1;
10347: pixelout<=1'b1;
10348: pixelout<=1'b1;
10349: pixelout<=1'b1;
10350: pixelout<=1'b1;
10351: pixelout<=1'b1;
10352: pixelout<=1'b1;
10353: pixelout<=1'b1;
10354: pixelout<=1'b1;
10355: pixelout<=1'b1;
10356: pixelout<=1'b1;
10357: pixelout<=1'b1;
10358: pixelout<=1'b1;
10359: pixelout<=1'b1;
10360: pixelout<=1'b1;
10361: pixelout<=1'b1;
10362: pixelout<=1'b1;
10363: pixelout<=1'b1;
10364: pixelout<=1'b1;
10365: pixelout<=1'b1;
10366: pixelout<=1'b1;
10367: pixelout<=1'b1;
10368: pixelout<=1'b1;
10369: pixelout<=1'b1;
10370: pixelout<=1'b1;
10371: pixelout<=1'b1;
10372: pixelout<=1'b1;
10373: pixelout<=1'b1;
10374: pixelout<=1'b1;
10375: pixelout<=1'b1;
10376: pixelout<=1'b1;
10377: pixelout<=1'b1;
10378: pixelout<=1'b1;
10379: pixelout<=1'b1;
10380: pixelout<=1'b1;
10381: pixelout<=1'b1;
10382: pixelout<=1'b1;
10383: pixelout<=1'b1;
10384: pixelout<=1'b1;
10385: pixelout<=1'b1;
10386: pixelout<=1'b1;
10387: pixelout<=1'b1;
10388: pixelout<=1'b1;
10389: pixelout<=1'b1;
10390: pixelout<=1'b1;
10391: pixelout<=1'b1;
10392: pixelout<=1'b1;
10393: pixelout<=1'b1;
10394: pixelout<=1'b1;
10395: pixelout<=1'b1;
10396: pixelout<=1'b1;
10397: pixelout<=1'b1;
10398: pixelout<=1'b1;
10399: pixelout<=1'b1;
10400: pixelout<=1'b1;
10401: pixelout<=1'b1;
10402: pixelout<=1'b1;
10403: pixelout<=1'b1;
10404: pixelout<=1'b1;
10405: pixelout<=1'b1;
10406: pixelout<=1'b1;
10407: pixelout<=1'b1;
10408: pixelout<=1'b1;
10409: pixelout<=1'b1;
10410: pixelout<=1'b1;
10411: pixelout<=1'b1;
10412: pixelout<=1'b1;
10413: pixelout<=1'b1;
10414: pixelout<=1'b1;
10415: pixelout<=1'b1;
10416: pixelout<=1'b1;
10417: pixelout<=1'b1;
10418: pixelout<=1'b1;
10419: pixelout<=1'b1;
10420: pixelout<=1'b1;
10421: pixelout<=1'b1;
10422: pixelout<=1'b1;
10423: pixelout<=1'b1;
10424: pixelout<=1'b1;
10425: pixelout<=1'b1;
10426: pixelout<=1'b1;
10427: pixelout<=1'b1;
10428: pixelout<=1'b1;
10429: pixelout<=1'b1;
10430: pixelout<=1'b1;
10431: pixelout<=1'b1;
10432: pixelout<=1'b1;
10433: pixelout<=1'b1;
10434: pixelout<=1'b1;
10435: pixelout<=1'b1;
10436: pixelout<=1'b1;
10437: pixelout<=1'b1;
10438: pixelout<=1'b1;
10439: pixelout<=1'b1;
10440: pixelout<=1'b1;
10441: pixelout<=1'b1;
10442: pixelout<=1'b1;
10443: pixelout<=1'b1;
10444: pixelout<=1'b1;
10445: pixelout<=1'b1;
10446: pixelout<=1'b1;
10447: pixelout<=1'b1;
10448: pixelout<=1'b1;
10449: pixelout<=1'b1;
10450: pixelout<=1'b1;
10451: pixelout<=1'b1;
10452: pixelout<=1'b1;
10453: pixelout<=1'b1;
10454: pixelout<=1'b1;
10455: pixelout<=1'b1;
10456: pixelout<=1'b1;
10457: pixelout<=1'b1;
10458: pixelout<=1'b1;
10459: pixelout<=1'b1;
10460: pixelout<=1'b1;
10461: pixelout<=1'b1;
10462: pixelout<=1'b1;
10463: pixelout<=1'b1;
10464: pixelout<=1'b1;
10465: pixelout<=1'b1;
10466: pixelout<=1'b1;
10467: pixelout<=1'b1;
10468: pixelout<=1'b1;
10469: pixelout<=1'b1;
10470: pixelout<=1'b1;
10471: pixelout<=1'b1;
10472: pixelout<=1'b1;
10473: pixelout<=1'b1;
10474: pixelout<=1'b1;
10475: pixelout<=1'b1;
10476: pixelout<=1'b1;
10477: pixelout<=1'b1;
10478: pixelout<=1'b1;
10479: pixelout<=1'b1;
10480: pixelout<=1'b1;
10481: pixelout<=1'b1;
10482: pixelout<=1'b1;
10483: pixelout<=1'b1;
10484: pixelout<=1'b1;
10485: pixelout<=1'b1;
10486: pixelout<=1'b1;
10487: pixelout<=1'b1;
10488: pixelout<=1'b1;
10489: pixelout<=1'b1;
10490: pixelout<=1'b1;
10491: pixelout<=1'b1;
10492: pixelout<=1'b1;
10493: pixelout<=1'b1;
10494: pixelout<=1'b1;
10495: pixelout<=1'b1;
10496: pixelout<=1'b1;
10497: pixelout<=1'b1;
10498: pixelout<=1'b1;
10499: pixelout<=1'b1;
10500: pixelout<=1'b1;
10501: pixelout<=1'b1;
10502: pixelout<=1'b1;
10503: pixelout<=1'b1;
10504: pixelout<=1'b1;
10505: pixelout<=1'b1;
10506: pixelout<=1'b1;
10507: pixelout<=1'b1;
10508: pixelout<=1'b1;
10509: pixelout<=1'b1;
10510: pixelout<=1'b1;
10511: pixelout<=1'b1;
10512: pixelout<=1'b1;
10513: pixelout<=1'b1;
10514: pixelout<=1'b1;
10515: pixelout<=1'b1;
10516: pixelout<=1'b1;
10517: pixelout<=1'b1;
10518: pixelout<=1'b1;
10519: pixelout<=1'b1;
10520: pixelout<=1'b1;
10521: pixelout<=1'b1;
10522: pixelout<=1'b1;
10523: pixelout<=1'b1;
10524: pixelout<=1'b1;
10525: pixelout<=1'b1;
10526: pixelout<=1'b1;
10527: pixelout<=1'b1;
10528: pixelout<=1'b1;
10529: pixelout<=1'b1;
10530: pixelout<=1'b1;
10531: pixelout<=1'b1;
10532: pixelout<=1'b1;
10533: pixelout<=1'b1;
10534: pixelout<=1'b1;
10535: pixelout<=1'b1;
10536: pixelout<=1'b1;
10537: pixelout<=1'b1;
10538: pixelout<=1'b1;
10539: pixelout<=1'b1;
10540: pixelout<=1'b1;
10541: pixelout<=1'b1;
10542: pixelout<=1'b1;
10543: pixelout<=1'b1;
10544: pixelout<=1'b1;
10545: pixelout<=1'b1;
10546: pixelout<=1'b1;
10547: pixelout<=1'b1;
10548: pixelout<=1'b1;
10549: pixelout<=1'b1;
10550: pixelout<=1'b1;
10551: pixelout<=1'b1;
10552: pixelout<=1'b1;
10553: pixelout<=1'b1;
10554: pixelout<=1'b1;
10555: pixelout<=1'b1;
10556: pixelout<=1'b1;
10557: pixelout<=1'b1;
10558: pixelout<=1'b1;
10559: pixelout<=1'b1;
10560: pixelout<=1'b1;
10561: pixelout<=1'b1;
10562: pixelout<=1'b1;
10563: pixelout<=1'b1;
10564: pixelout<=1'b1;
10565: pixelout<=1'b1;
10566: pixelout<=1'b1;
10567: pixelout<=1'b1;
10568: pixelout<=1'b1;
10569: pixelout<=1'b1;
10570: pixelout<=1'b1;
10571: pixelout<=1'b1;
10572: pixelout<=1'b1;
10573: pixelout<=1'b1;
10574: pixelout<=1'b1;
10575: pixelout<=1'b1;
10576: pixelout<=1'b1;
10577: pixelout<=1'b1;
10578: pixelout<=1'b1;
10579: pixelout<=1'b1;
10580: pixelout<=1'b1;
10581: pixelout<=1'b1;
10582: pixelout<=1'b1;
10583: pixelout<=1'b1;
10584: pixelout<=1'b1;
10585: pixelout<=1'b1;
10586: pixelout<=1'b1;
10587: pixelout<=1'b1;
10588: pixelout<=1'b1;
10589: pixelout<=1'b1;
10590: pixelout<=1'b1;
10591: pixelout<=1'b1;
10592: pixelout<=1'b1;
10593: pixelout<=1'b1;
10594: pixelout<=1'b1;
10595: pixelout<=1'b1;
10596: pixelout<=1'b1;
10597: pixelout<=1'b1;
10598: pixelout<=1'b1;
10599: pixelout<=1'b1;
10600: pixelout<=1'b1;
10601: pixelout<=1'b1;
10602: pixelout<=1'b1;
10603: pixelout<=1'b1;
10604: pixelout<=1'b1;
10605: pixelout<=1'b1;
10606: pixelout<=1'b1;
10607: pixelout<=1'b1;
10608: pixelout<=1'b1;
10609: pixelout<=1'b1;
10610: pixelout<=1'b1;
10611: pixelout<=1'b1;
10612: pixelout<=1'b1;
10613: pixelout<=1'b1;
10614: pixelout<=1'b1;
10615: pixelout<=1'b1;
10616: pixelout<=1'b1;
10617: pixelout<=1'b1;
10618: pixelout<=1'b1;
10619: pixelout<=1'b1;
10620: pixelout<=1'b1;
10621: pixelout<=1'b1;
10622: pixelout<=1'b1;
10623: pixelout<=1'b1;
10624: pixelout<=1'b1;
10625: pixelout<=1'b1;
10626: pixelout<=1'b1;
10627: pixelout<=1'b1;
10628: pixelout<=1'b1;
10629: pixelout<=1'b1;
10630: pixelout<=1'b1;
10631: pixelout<=1'b1;
10632: pixelout<=1'b1;
10633: pixelout<=1'b1;
10634: pixelout<=1'b1;
10635: pixelout<=1'b1;
10636: pixelout<=1'b1;
10637: pixelout<=1'b1;
10638: pixelout<=1'b1;
10639: pixelout<=1'b1;
10640: pixelout<=1'b1;
10641: pixelout<=1'b1;
10642: pixelout<=1'b1;
10643: pixelout<=1'b1;
10644: pixelout<=1'b1;
10645: pixelout<=1'b1;
10646: pixelout<=1'b1;
10647: pixelout<=1'b1;
10648: pixelout<=1'b1;
10649: pixelout<=1'b1;
10650: pixelout<=1'b1;
10651: pixelout<=1'b1;
10652: pixelout<=1'b1;
10653: pixelout<=1'b1;
10654: pixelout<=1'b1;
10655: pixelout<=1'b1;
10656: pixelout<=1'b1;
10657: pixelout<=1'b1;
10658: pixelout<=1'b1;
10659: pixelout<=1'b1;
10660: pixelout<=1'b1;
10661: pixelout<=1'b1;
10662: pixelout<=1'b1;
10663: pixelout<=1'b1;
10664: pixelout<=1'b1;
10665: pixelout<=1'b1;
10666: pixelout<=1'b1;
10667: pixelout<=1'b1;
10668: pixelout<=1'b1;
10669: pixelout<=1'b1;
10670: pixelout<=1'b1;
10671: pixelout<=1'b1;
10672: pixelout<=1'b1;
10673: pixelout<=1'b1;
10674: pixelout<=1'b1;
10675: pixelout<=1'b1;
10676: pixelout<=1'b1;
10677: pixelout<=1'b1;
10678: pixelout<=1'b1;
10679: pixelout<=1'b1;
10680: pixelout<=1'b1;
10681: pixelout<=1'b1;
10682: pixelout<=1'b1;
10683: pixelout<=1'b1;
10684: pixelout<=1'b1;
10685: pixelout<=1'b1;
10686: pixelout<=1'b1;
10687: pixelout<=1'b1;
10688: pixelout<=1'b1;
10689: pixelout<=1'b1;
10690: pixelout<=1'b1;
10691: pixelout<=1'b1;
10692: pixelout<=1'b1;
10693: pixelout<=1'b1;
10694: pixelout<=1'b1;
10695: pixelout<=1'b1;
10696: pixelout<=1'b1;
10697: pixelout<=1'b1;
10698: pixelout<=1'b1;
10699: pixelout<=1'b1;
10700: pixelout<=1'b1;
10701: pixelout<=1'b1;
10702: pixelout<=1'b1;
10703: pixelout<=1'b1;
10704: pixelout<=1'b1;
10705: pixelout<=1'b1;
10706: pixelout<=1'b1;
10707: pixelout<=1'b1;
10708: pixelout<=1'b1;
10709: pixelout<=1'b1;
10710: pixelout<=1'b1;
10711: pixelout<=1'b1;
10712: pixelout<=1'b1;
10713: pixelout<=1'b1;
10714: pixelout<=1'b1;
10715: pixelout<=1'b1;
10716: pixelout<=1'b1;
10717: pixelout<=1'b1;
10718: pixelout<=1'b1;
10719: pixelout<=1'b1;
10720: pixelout<=1'b1;
10721: pixelout<=1'b1;
10722: pixelout<=1'b1;
10723: pixelout<=1'b1;
10724: pixelout<=1'b1;
10725: pixelout<=1'b1;
10726: pixelout<=1'b1;
10727: pixelout<=1'b1;
10728: pixelout<=1'b1;
10729: pixelout<=1'b1;
10730: pixelout<=1'b1;
10731: pixelout<=1'b1;
10732: pixelout<=1'b1;
10733: pixelout<=1'b1;
10734: pixelout<=1'b1;
10735: pixelout<=1'b1;
10736: pixelout<=1'b1;
10737: pixelout<=1'b1;
10738: pixelout<=1'b1;
10739: pixelout<=1'b1;
10740: pixelout<=1'b1;
10741: pixelout<=1'b1;
10742: pixelout<=1'b1;
10743: pixelout<=1'b1;
10744: pixelout<=1'b1;
10745: pixelout<=1'b1;
10746: pixelout<=1'b1;
10747: pixelout<=1'b1;
10748: pixelout<=1'b1;
10749: pixelout<=1'b1;
10750: pixelout<=1'b1;
10751: pixelout<=1'b1;
10752: pixelout<=1'b1;
10753: pixelout<=1'b1;
10754: pixelout<=1'b1;
10755: pixelout<=1'b1;
10756: pixelout<=1'b1;
10757: pixelout<=1'b1;
10758: pixelout<=1'b1;
10759: pixelout<=1'b1;
10760: pixelout<=1'b1;
10761: pixelout<=1'b1;
10762: pixelout<=1'b1;
10763: pixelout<=1'b1;
10764: pixelout<=1'b1;
10765: pixelout<=1'b1;
10766: pixelout<=1'b1;
10767: pixelout<=1'b1;
10768: pixelout<=1'b1;
10769: pixelout<=1'b1;
10770: pixelout<=1'b1;
10771: pixelout<=1'b1;
10772: pixelout<=1'b1;
10773: pixelout<=1'b1;
10774: pixelout<=1'b1;
10775: pixelout<=1'b1;
10776: pixelout<=1'b1;
10777: pixelout<=1'b1;
10778: pixelout<=1'b1;
10779: pixelout<=1'b1;
10780: pixelout<=1'b1;
10781: pixelout<=1'b1;
10782: pixelout<=1'b1;
10783: pixelout<=1'b1;
10784: pixelout<=1'b1;
10785: pixelout<=1'b1;
10786: pixelout<=1'b1;
10787: pixelout<=1'b1;
10788: pixelout<=1'b1;
10789: pixelout<=1'b1;
10790: pixelout<=1'b1;
10791: pixelout<=1'b1;
10792: pixelout<=1'b1;
10793: pixelout<=1'b1;
10794: pixelout<=1'b1;
10795: pixelout<=1'b1;
10796: pixelout<=1'b1;
10797: pixelout<=1'b1;
10798: pixelout<=1'b1;
10799: pixelout<=1'b1;
10800: pixelout<=1'b1;
10801: pixelout<=1'b1;
10802: pixelout<=1'b1;
10803: pixelout<=1'b1;
10804: pixelout<=1'b1;
10805: pixelout<=1'b1;
10806: pixelout<=1'b1;
10807: pixelout<=1'b1;
10808: pixelout<=1'b1;
10809: pixelout<=1'b1;
10810: pixelout<=1'b1;
10811: pixelout<=1'b1;
10812: pixelout<=1'b1;
10813: pixelout<=1'b1;
10814: pixelout<=1'b1;
10815: pixelout<=1'b1;
10816: pixelout<=1'b1;
10817: pixelout<=1'b1;
10818: pixelout<=1'b1;
10819: pixelout<=1'b1;
10820: pixelout<=1'b1;
10821: pixelout<=1'b1;
10822: pixelout<=1'b1;
10823: pixelout<=1'b1;
10824: pixelout<=1'b1;
10825: pixelout<=1'b1;
10826: pixelout<=1'b1;
10827: pixelout<=1'b1;
10828: pixelout<=1'b1;
10829: pixelout<=1'b1;
10830: pixelout<=1'b1;
10831: pixelout<=1'b1;
10832: pixelout<=1'b1;
10833: pixelout<=1'b1;
10834: pixelout<=1'b1;
10835: pixelout<=1'b1;
10836: pixelout<=1'b1;
10837: pixelout<=1'b1;
10838: pixelout<=1'b1;
10839: pixelout<=1'b1;
10840: pixelout<=1'b1;
10841: pixelout<=1'b1;
10842: pixelout<=1'b1;
10843: pixelout<=1'b1;
10844: pixelout<=1'b1;
10845: pixelout<=1'b1;
10846: pixelout<=1'b1;
10847: pixelout<=1'b1;
10848: pixelout<=1'b1;
10849: pixelout<=1'b1;
10850: pixelout<=1'b1;
10851: pixelout<=1'b1;
10852: pixelout<=1'b1;
10853: pixelout<=1'b1;
10854: pixelout<=1'b1;
10855: pixelout<=1'b1;
10856: pixelout<=1'b1;
10857: pixelout<=1'b1;
10858: pixelout<=1'b1;
10859: pixelout<=1'b1;
10860: pixelout<=1'b1;
10861: pixelout<=1'b1;
10862: pixelout<=1'b1;
10863: pixelout<=1'b1;
10864: pixelout<=1'b1;
10865: pixelout<=1'b1;
10866: pixelout<=1'b1;
10867: pixelout<=1'b1;
10868: pixelout<=1'b1;
10869: pixelout<=1'b1;
10870: pixelout<=1'b1;
10871: pixelout<=1'b1;
10872: pixelout<=1'b1;
10873: pixelout<=1'b1;
10874: pixelout<=1'b1;
10875: pixelout<=1'b1;
10876: pixelout<=1'b1;
10877: pixelout<=1'b1;
10878: pixelout<=1'b1;
10879: pixelout<=1'b1;
10880: pixelout<=1'b1;
10881: pixelout<=1'b1;
10882: pixelout<=1'b1;
10883: pixelout<=1'b1;
10884: pixelout<=1'b1;
10885: pixelout<=1'b1;
10886: pixelout<=1'b1;
10887: pixelout<=1'b1;
10888: pixelout<=1'b1;
10889: pixelout<=1'b1;
10890: pixelout<=1'b1;
10891: pixelout<=1'b1;
10892: pixelout<=1'b1;
10893: pixelout<=1'b1;
10894: pixelout<=1'b1;
10895: pixelout<=1'b1;
10896: pixelout<=1'b1;
10897: pixelout<=1'b1;
10898: pixelout<=1'b1;
10899: pixelout<=1'b1;
10900: pixelout<=1'b1;
10901: pixelout<=1'b1;
10902: pixelout<=1'b1;
10903: pixelout<=1'b1;
10904: pixelout<=1'b1;
10905: pixelout<=1'b1;
10906: pixelout<=1'b1;
10907: pixelout<=1'b1;
10908: pixelout<=1'b1;
10909: pixelout<=1'b1;
10910: pixelout<=1'b1;
10911: pixelout<=1'b1;
10912: pixelout<=1'b1;
10913: pixelout<=1'b1;
10914: pixelout<=1'b1;
10915: pixelout<=1'b1;
10916: pixelout<=1'b1;
10917: pixelout<=1'b1;
10918: pixelout<=1'b1;
10919: pixelout<=1'b1;
10920: pixelout<=1'b1;
10921: pixelout<=1'b1;
10922: pixelout<=1'b1;
10923: pixelout<=1'b1;
10924: pixelout<=1'b1;
10925: pixelout<=1'b1;
10926: pixelout<=1'b1;
10927: pixelout<=1'b1;
10928: pixelout<=1'b1;
10929: pixelout<=1'b1;
10930: pixelout<=1'b1;
10931: pixelout<=1'b1;
10932: pixelout<=1'b1;
10933: pixelout<=1'b1;
10934: pixelout<=1'b1;
10935: pixelout<=1'b1;
10936: pixelout<=1'b1;
10937: pixelout<=1'b1;
10938: pixelout<=1'b1;
10939: pixelout<=1'b1;
10940: pixelout<=1'b1;
10941: pixelout<=1'b1;
10942: pixelout<=1'b1;
10943: pixelout<=1'b1;
10944: pixelout<=1'b1;
10945: pixelout<=1'b1;
10946: pixelout<=1'b1;
10947: pixelout<=1'b1;
10948: pixelout<=1'b1;
10949: pixelout<=1'b1;
10950: pixelout<=1'b1;
10951: pixelout<=1'b1;
10952: pixelout<=1'b1;
10953: pixelout<=1'b1;
10954: pixelout<=1'b1;
10955: pixelout<=1'b1;
10956: pixelout<=1'b1;
10957: pixelout<=1'b1;
10958: pixelout<=1'b1;
10959: pixelout<=1'b1;
10960: pixelout<=1'b1;
10961: pixelout<=1'b1;
10962: pixelout<=1'b1;
10963: pixelout<=1'b1;
10964: pixelout<=1'b1;
10965: pixelout<=1'b1;
10966: pixelout<=1'b1;
10967: pixelout<=1'b1;
10968: pixelout<=1'b1;
10969: pixelout<=1'b1;
10970: pixelout<=1'b1;
10971: pixelout<=1'b1;
10972: pixelout<=1'b1;
10973: pixelout<=1'b1;
10974: pixelout<=1'b1;
10975: pixelout<=1'b1;
10976: pixelout<=1'b1;
10977: pixelout<=1'b1;
10978: pixelout<=1'b1;
10979: pixelout<=1'b1;
10980: pixelout<=1'b1;
10981: pixelout<=1'b1;
10982: pixelout<=1'b1;
10983: pixelout<=1'b1;
10984: pixelout<=1'b1;
10985: pixelout<=1'b1;
10986: pixelout<=1'b1;
10987: pixelout<=1'b1;
10988: pixelout<=1'b1;
10989: pixelout<=1'b1;
10990: pixelout<=1'b1;
10991: pixelout<=1'b1;
10992: pixelout<=1'b1;
10993: pixelout<=1'b1;
10994: pixelout<=1'b1;
10995: pixelout<=1'b1;
10996: pixelout<=1'b1;
10997: pixelout<=1'b1;
10998: pixelout<=1'b1;
10999: pixelout<=1'b1;
11000: pixelout<=1'b1;
11001: pixelout<=1'b1;
11002: pixelout<=1'b1;
11003: pixelout<=1'b1;
11004: pixelout<=1'b1;
11005: pixelout<=1'b1;
11006: pixelout<=1'b1;
11007: pixelout<=1'b1;
11008: pixelout<=1'b1;
11009: pixelout<=1'b1;
11010: pixelout<=1'b1;
11011: pixelout<=1'b1;
11012: pixelout<=1'b1;
11013: pixelout<=1'b1;
11014: pixelout<=1'b1;
11015: pixelout<=1'b1;
11016: pixelout<=1'b1;
11017: pixelout<=1'b1;
11018: pixelout<=1'b1;
11019: pixelout<=1'b1;
11020: pixelout<=1'b1;
11021: pixelout<=1'b1;
11022: pixelout<=1'b1;
11023: pixelout<=1'b1;
11024: pixelout<=1'b1;
11025: pixelout<=1'b1;
11026: pixelout<=1'b1;
11027: pixelout<=1'b1;
11028: pixelout<=1'b1;
11029: pixelout<=1'b1;
11030: pixelout<=1'b1;
11031: pixelout<=1'b1;
11032: pixelout<=1'b1;
11033: pixelout<=1'b1;
11034: pixelout<=1'b1;
11035: pixelout<=1'b1;
11036: pixelout<=1'b1;
11037: pixelout<=1'b1;
11038: pixelout<=1'b1;
11039: pixelout<=1'b1;
11040: pixelout<=1'b1;
11041: pixelout<=1'b1;
11042: pixelout<=1'b1;
11043: pixelout<=1'b1;
11044: pixelout<=1'b1;
11045: pixelout<=1'b1;
11046: pixelout<=1'b1;
11047: pixelout<=1'b1;
11048: pixelout<=1'b1;
11049: pixelout<=1'b1;
11050: pixelout<=1'b1;
11051: pixelout<=1'b1;
11052: pixelout<=1'b1;
11053: pixelout<=1'b1;
11054: pixelout<=1'b1;
11055: pixelout<=1'b1;
11056: pixelout<=1'b1;
11057: pixelout<=1'b1;
11058: pixelout<=1'b1;
11059: pixelout<=1'b1;
11060: pixelout<=1'b1;
11061: pixelout<=1'b1;
11062: pixelout<=1'b1;
11063: pixelout<=1'b1;
11064: pixelout<=1'b1;
11065: pixelout<=1'b1;
11066: pixelout<=1'b1;
11067: pixelout<=1'b1;
11068: pixelout<=1'b1;
11069: pixelout<=1'b1;
11070: pixelout<=1'b1;
11071: pixelout<=1'b1;
11072: pixelout<=1'b1;
11073: pixelout<=1'b1;
11074: pixelout<=1'b1;
11075: pixelout<=1'b1;
11076: pixelout<=1'b1;
11077: pixelout<=1'b1;
11078: pixelout<=1'b1;
11079: pixelout<=1'b1;
11080: pixelout<=1'b1;
11081: pixelout<=1'b1;
11082: pixelout<=1'b1;
11083: pixelout<=1'b1;
11084: pixelout<=1'b1;
11085: pixelout<=1'b1;
11086: pixelout<=1'b1;
11087: pixelout<=1'b1;
11088: pixelout<=1'b1;
11089: pixelout<=1'b1;
11090: pixelout<=1'b1;
11091: pixelout<=1'b1;
11092: pixelout<=1'b1;
11093: pixelout<=1'b1;
11094: pixelout<=1'b1;
11095: pixelout<=1'b1;
11096: pixelout<=1'b1;
11097: pixelout<=1'b1;
11098: pixelout<=1'b1;
11099: pixelout<=1'b1;
11100: pixelout<=1'b1;
11101: pixelout<=1'b1;
11102: pixelout<=1'b1;
11103: pixelout<=1'b1;
11104: pixelout<=1'b1;
11105: pixelout<=1'b1;
11106: pixelout<=1'b1;
11107: pixelout<=1'b1;
11108: pixelout<=1'b1;
11109: pixelout<=1'b1;
11110: pixelout<=1'b1;
11111: pixelout<=1'b1;
11112: pixelout<=1'b1;
11113: pixelout<=1'b1;
11114: pixelout<=1'b1;
11115: pixelout<=1'b1;
11116: pixelout<=1'b1;
11117: pixelout<=1'b1;
11118: pixelout<=1'b1;
11119: pixelout<=1'b1;
11120: pixelout<=1'b1;
11121: pixelout<=1'b1;
11122: pixelout<=1'b1;
11123: pixelout<=1'b1;
11124: pixelout<=1'b1;
11125: pixelout<=1'b1;
11126: pixelout<=1'b1;
11127: pixelout<=1'b1;
11128: pixelout<=1'b1;
11129: pixelout<=1'b1;
11130: pixelout<=1'b1;
11131: pixelout<=1'b1;
11132: pixelout<=1'b1;
11133: pixelout<=1'b1;
11134: pixelout<=1'b1;
11135: pixelout<=1'b1;
11136: pixelout<=1'b1;
11137: pixelout<=1'b1;
11138: pixelout<=1'b1;
11139: pixelout<=1'b1;
11140: pixelout<=1'b1;
11141: pixelout<=1'b1;
11142: pixelout<=1'b1;
11143: pixelout<=1'b1;
11144: pixelout<=1'b1;
11145: pixelout<=1'b1;
11146: pixelout<=1'b1;
11147: pixelout<=1'b1;
11148: pixelout<=1'b1;
11149: pixelout<=1'b1;
11150: pixelout<=1'b1;
11151: pixelout<=1'b1;
11152: pixelout<=1'b1;
11153: pixelout<=1'b1;
11154: pixelout<=1'b1;
11155: pixelout<=1'b1;
11156: pixelout<=1'b1;
11157: pixelout<=1'b1;
11158: pixelout<=1'b1;
11159: pixelout<=1'b1;
11160: pixelout<=1'b1;
11161: pixelout<=1'b1;
11162: pixelout<=1'b1;
11163: pixelout<=1'b1;
11164: pixelout<=1'b1;
11165: pixelout<=1'b1;
11166: pixelout<=1'b1;
11167: pixelout<=1'b1;
11168: pixelout<=1'b1;
11169: pixelout<=1'b1;
11170: pixelout<=1'b1;
11171: pixelout<=1'b1;
11172: pixelout<=1'b1;
11173: pixelout<=1'b1;
11174: pixelout<=1'b1;
11175: pixelout<=1'b1;
11176: pixelout<=1'b1;
11177: pixelout<=1'b1;
11178: pixelout<=1'b1;
11179: pixelout<=1'b1;
11180: pixelout<=1'b1;
11181: pixelout<=1'b1;
11182: pixelout<=1'b1;
11183: pixelout<=1'b1;
11184: pixelout<=1'b1;
11185: pixelout<=1'b1;
11186: pixelout<=1'b1;
11187: pixelout<=1'b1;
11188: pixelout<=1'b1;
11189: pixelout<=1'b1;
11190: pixelout<=1'b1;
11191: pixelout<=1'b1;
11192: pixelout<=1'b1;
11193: pixelout<=1'b1;
11194: pixelout<=1'b1;
11195: pixelout<=1'b1;
11196: pixelout<=1'b1;
11197: pixelout<=1'b1;
11198: pixelout<=1'b1;
11199: pixelout<=1'b1;
11200: pixelout<=1'b1;
11201: pixelout<=1'b1;
11202: pixelout<=1'b1;
11203: pixelout<=1'b1;
11204: pixelout<=1'b1;
11205: pixelout<=1'b1;
11206: pixelout<=1'b1;
11207: pixelout<=1'b1;
11208: pixelout<=1'b1;
11209: pixelout<=1'b1;
11210: pixelout<=1'b1;
11211: pixelout<=1'b1;
11212: pixelout<=1'b1;
11213: pixelout<=1'b1;
11214: pixelout<=1'b1;
11215: pixelout<=1'b1;
11216: pixelout<=1'b1;
11217: pixelout<=1'b1;
11218: pixelout<=1'b1;
11219: pixelout<=1'b1;
11220: pixelout<=1'b1;
11221: pixelout<=1'b1;
11222: pixelout<=1'b1;
11223: pixelout<=1'b1;
11224: pixelout<=1'b1;
11225: pixelout<=1'b1;
11226: pixelout<=1'b1;
11227: pixelout<=1'b1;
11228: pixelout<=1'b1;
11229: pixelout<=1'b1;
11230: pixelout<=1'b1;
11231: pixelout<=1'b1;
11232: pixelout<=1'b1;
11233: pixelout<=1'b1;
11234: pixelout<=1'b1;
11235: pixelout<=1'b1;
11236: pixelout<=1'b1;
11237: pixelout<=1'b1;
11238: pixelout<=1'b1;
11239: pixelout<=1'b1;
11240: pixelout<=1'b1;
11241: pixelout<=1'b1;
11242: pixelout<=1'b1;
11243: pixelout<=1'b1;
11244: pixelout<=1'b1;
11245: pixelout<=1'b1;
11246: pixelout<=1'b1;
11247: pixelout<=1'b1;
11248: pixelout<=1'b1;
11249: pixelout<=1'b1;
11250: pixelout<=1'b1;
11251: pixelout<=1'b1;
11252: pixelout<=1'b1;
11253: pixelout<=1'b1;
11254: pixelout<=1'b1;
11255: pixelout<=1'b1;
11256: pixelout<=1'b1;
11257: pixelout<=1'b1;
11258: pixelout<=1'b1;
11259: pixelout<=1'b1;
11260: pixelout<=1'b1;
11261: pixelout<=1'b1;
11262: pixelout<=1'b1;
11263: pixelout<=1'b1;
11264: pixelout<=1'b1;
11265: pixelout<=1'b1;
11266: pixelout<=1'b1;
11267: pixelout<=1'b1;
11268: pixelout<=1'b1;
11269: pixelout<=1'b1;
11270: pixelout<=1'b1;
11271: pixelout<=1'b1;
11272: pixelout<=1'b1;
11273: pixelout<=1'b1;
11274: pixelout<=1'b1;
11275: pixelout<=1'b1;
11276: pixelout<=1'b1;
11277: pixelout<=1'b1;
11278: pixelout<=1'b1;
11279: pixelout<=1'b1;
11280: pixelout<=1'b1;
11281: pixelout<=1'b1;
11282: pixelout<=1'b1;
11283: pixelout<=1'b1;
11284: pixelout<=1'b1;
11285: pixelout<=1'b1;
11286: pixelout<=1'b1;
11287: pixelout<=1'b1;
11288: pixelout<=1'b1;
11289: pixelout<=1'b1;
11290: pixelout<=1'b1;
11291: pixelout<=1'b1;
11292: pixelout<=1'b1;
11293: pixelout<=1'b1;
11294: pixelout<=1'b1;
11295: pixelout<=1'b1;
11296: pixelout<=1'b1;
11297: pixelout<=1'b1;
11298: pixelout<=1'b1;
11299: pixelout<=1'b1;
11300: pixelout<=1'b1;
11301: pixelout<=1'b1;
11302: pixelout<=1'b1;
11303: pixelout<=1'b1;
11304: pixelout<=1'b1;
11305: pixelout<=1'b1;
11306: pixelout<=1'b1;
11307: pixelout<=1'b1;
11308: pixelout<=1'b1;
11309: pixelout<=1'b1;
11310: pixelout<=1'b1;
11311: pixelout<=1'b1;
11312: pixelout<=1'b1;
11313: pixelout<=1'b1;
11314: pixelout<=1'b1;
11315: pixelout<=1'b1;
11316: pixelout<=1'b1;
11317: pixelout<=1'b1;
11318: pixelout<=1'b1;
11319: pixelout<=1'b1;
11320: pixelout<=1'b1;
11321: pixelout<=1'b1;
11322: pixelout<=1'b1;
11323: pixelout<=1'b1;
11324: pixelout<=1'b1;
11325: pixelout<=1'b1;
11326: pixelout<=1'b1;
11327: pixelout<=1'b1;
11328: pixelout<=1'b1;
11329: pixelout<=1'b1;
11330: pixelout<=1'b1;
11331: pixelout<=1'b1;
11332: pixelout<=1'b1;
11333: pixelout<=1'b1;
11334: pixelout<=1'b1;
11335: pixelout<=1'b1;
11336: pixelout<=1'b1;
11337: pixelout<=1'b1;
11338: pixelout<=1'b1;
11339: pixelout<=1'b1;
11340: pixelout<=1'b1;
11341: pixelout<=1'b1;
11342: pixelout<=1'b1;
11343: pixelout<=1'b1;
11344: pixelout<=1'b1;
11345: pixelout<=1'b1;
11346: pixelout<=1'b1;
11347: pixelout<=1'b1;
11348: pixelout<=1'b1;
11349: pixelout<=1'b1;
11350: pixelout<=1'b1;
11351: pixelout<=1'b1;
11352: pixelout<=1'b1;
11353: pixelout<=1'b1;
11354: pixelout<=1'b1;
11355: pixelout<=1'b1;
11356: pixelout<=1'b1;
11357: pixelout<=1'b1;
11358: pixelout<=1'b1;
11359: pixelout<=1'b1;
11360: pixelout<=1'b1;
11361: pixelout<=1'b1;
11362: pixelout<=1'b1;
11363: pixelout<=1'b1;
11364: pixelout<=1'b1;
11365: pixelout<=1'b1;
11366: pixelout<=1'b1;
11367: pixelout<=1'b1;
11368: pixelout<=1'b1;
11369: pixelout<=1'b1;
11370: pixelout<=1'b1;
11371: pixelout<=1'b1;
11372: pixelout<=1'b1;
11373: pixelout<=1'b1;
11374: pixelout<=1'b1;
11375: pixelout<=1'b1;
11376: pixelout<=1'b1;
11377: pixelout<=1'b1;
11378: pixelout<=1'b1;
11379: pixelout<=1'b1;
11380: pixelout<=1'b1;
11381: pixelout<=1'b1;
11382: pixelout<=1'b1;
11383: pixelout<=1'b1;
11384: pixelout<=1'b1;
11385: pixelout<=1'b1;
11386: pixelout<=1'b1;
11387: pixelout<=1'b1;
11388: pixelout<=1'b1;
11389: pixelout<=1'b1;
11390: pixelout<=1'b1;
11391: pixelout<=1'b1;
11392: pixelout<=1'b1;
11393: pixelout<=1'b1;
11394: pixelout<=1'b1;
11395: pixelout<=1'b1;
11396: pixelout<=1'b1;
11397: pixelout<=1'b1;
11398: pixelout<=1'b1;
11399: pixelout<=1'b1;
11400: pixelout<=1'b1;
11401: pixelout<=1'b1;
11402: pixelout<=1'b1;
11403: pixelout<=1'b1;
11404: pixelout<=1'b1;
11405: pixelout<=1'b1;
11406: pixelout<=1'b1;
11407: pixelout<=1'b1;
11408: pixelout<=1'b1;
11409: pixelout<=1'b1;
11410: pixelout<=1'b1;
11411: pixelout<=1'b1;
11412: pixelout<=1'b1;
11413: pixelout<=1'b1;
11414: pixelout<=1'b1;
11415: pixelout<=1'b1;
11416: pixelout<=1'b1;
11417: pixelout<=1'b1;
11418: pixelout<=1'b1;
11419: pixelout<=1'b1;
11420: pixelout<=1'b1;
11421: pixelout<=1'b1;
11422: pixelout<=1'b1;
11423: pixelout<=1'b1;
11424: pixelout<=1'b1;
11425: pixelout<=1'b1;
11426: pixelout<=1'b1;
11427: pixelout<=1'b1;
11428: pixelout<=1'b1;
11429: pixelout<=1'b1;
11430: pixelout<=1'b1;
11431: pixelout<=1'b1;
11432: pixelout<=1'b1;
11433: pixelout<=1'b1;
11434: pixelout<=1'b1;
11435: pixelout<=1'b1;
11436: pixelout<=1'b1;
11437: pixelout<=1'b1;
11438: pixelout<=1'b1;
11439: pixelout<=1'b1;
11440: pixelout<=1'b1;
11441: pixelout<=1'b1;
11442: pixelout<=1'b1;
11443: pixelout<=1'b1;
11444: pixelout<=1'b1;
11445: pixelout<=1'b1;
11446: pixelout<=1'b1;
11447: pixelout<=1'b1;
11448: pixelout<=1'b1;
11449: pixelout<=1'b1;
11450: pixelout<=1'b1;
11451: pixelout<=1'b1;
11452: pixelout<=1'b1;
11453: pixelout<=1'b1;
11454: pixelout<=1'b1;
11455: pixelout<=1'b1;
11456: pixelout<=1'b1;
11457: pixelout<=1'b1;
11458: pixelout<=1'b1;
11459: pixelout<=1'b1;
11460: pixelout<=1'b1;
11461: pixelout<=1'b1;
11462: pixelout<=1'b1;
11463: pixelout<=1'b1;
11464: pixelout<=1'b1;
11465: pixelout<=1'b1;
11466: pixelout<=1'b1;
11467: pixelout<=1'b1;
11468: pixelout<=1'b1;
11469: pixelout<=1'b1;
11470: pixelout<=1'b1;
11471: pixelout<=1'b1;
11472: pixelout<=1'b1;
11473: pixelout<=1'b1;
11474: pixelout<=1'b1;
11475: pixelout<=1'b1;
11476: pixelout<=1'b1;
11477: pixelout<=1'b1;
11478: pixelout<=1'b1;
11479: pixelout<=1'b1;
11480: pixelout<=1'b1;
11481: pixelout<=1'b1;
11482: pixelout<=1'b1;
11483: pixelout<=1'b1;
11484: pixelout<=1'b1;
11485: pixelout<=1'b1;
11486: pixelout<=1'b1;
11487: pixelout<=1'b1;
11488: pixelout<=1'b1;
11489: pixelout<=1'b1;
11490: pixelout<=1'b1;
11491: pixelout<=1'b1;
11492: pixelout<=1'b1;
11493: pixelout<=1'b1;
11494: pixelout<=1'b1;
11495: pixelout<=1'b1;
11496: pixelout<=1'b1;
11497: pixelout<=1'b1;
11498: pixelout<=1'b1;
11499: pixelout<=1'b1;
11500: pixelout<=1'b1;
11501: pixelout<=1'b1;
11502: pixelout<=1'b1;
11503: pixelout<=1'b1;
11504: pixelout<=1'b1;
11505: pixelout<=1'b1;
11506: pixelout<=1'b1;
11507: pixelout<=1'b1;
11508: pixelout<=1'b1;
11509: pixelout<=1'b1;
11510: pixelout<=1'b1;
11511: pixelout<=1'b1;
11512: pixelout<=1'b1;
11513: pixelout<=1'b1;
11514: pixelout<=1'b1;
11515: pixelout<=1'b1;
11516: pixelout<=1'b1;
11517: pixelout<=1'b1;
11518: pixelout<=1'b1;
11519: pixelout<=1'b1;
11520: pixelout<=1'b1;
11521: pixelout<=1'b1;
11522: pixelout<=1'b1;
11523: pixelout<=1'b1;
11524: pixelout<=1'b1;
11525: pixelout<=1'b1;
11526: pixelout<=1'b1;
11527: pixelout<=1'b1;
11528: pixelout<=1'b1;
11529: pixelout<=1'b1;
11530: pixelout<=1'b1;
11531: pixelout<=1'b1;
11532: pixelout<=1'b1;
11533: pixelout<=1'b1;
11534: pixelout<=1'b1;
11535: pixelout<=1'b1;
11536: pixelout<=1'b1;
11537: pixelout<=1'b1;
11538: pixelout<=1'b1;
11539: pixelout<=1'b1;
11540: pixelout<=1'b1;
11541: pixelout<=1'b1;
11542: pixelout<=1'b1;
11543: pixelout<=1'b1;
11544: pixelout<=1'b1;
11545: pixelout<=1'b1;
11546: pixelout<=1'b1;
11547: pixelout<=1'b1;
11548: pixelout<=1'b1;
11549: pixelout<=1'b1;
11550: pixelout<=1'b1;
11551: pixelout<=1'b1;
11552: pixelout<=1'b1;
11553: pixelout<=1'b1;
11554: pixelout<=1'b1;
11555: pixelout<=1'b1;
11556: pixelout<=1'b1;
11557: pixelout<=1'b1;
11558: pixelout<=1'b1;
11559: pixelout<=1'b1;
11560: pixelout<=1'b1;
11561: pixelout<=1'b1;
11562: pixelout<=1'b1;
11563: pixelout<=1'b1;
11564: pixelout<=1'b1;
11565: pixelout<=1'b1;
11566: pixelout<=1'b1;
11567: pixelout<=1'b1;
11568: pixelout<=1'b1;
11569: pixelout<=1'b1;
11570: pixelout<=1'b1;
11571: pixelout<=1'b1;
11572: pixelout<=1'b1;
11573: pixelout<=1'b1;
11574: pixelout<=1'b1;
11575: pixelout<=1'b1;
11576: pixelout<=1'b1;
11577: pixelout<=1'b1;
11578: pixelout<=1'b1;
11579: pixelout<=1'b1;
11580: pixelout<=1'b1;
11581: pixelout<=1'b1;
11582: pixelout<=1'b1;
11583: pixelout<=1'b1;
11584: pixelout<=1'b1;
11585: pixelout<=1'b1;
11586: pixelout<=1'b1;
11587: pixelout<=1'b1;
11588: pixelout<=1'b1;
11589: pixelout<=1'b1;
11590: pixelout<=1'b1;
11591: pixelout<=1'b1;
11592: pixelout<=1'b1;
11593: pixelout<=1'b1;
11594: pixelout<=1'b1;
11595: pixelout<=1'b1;
11596: pixelout<=1'b1;
11597: pixelout<=1'b1;
11598: pixelout<=1'b1;
11599: pixelout<=1'b1;
11600: pixelout<=1'b1;
11601: pixelout<=1'b1;
11602: pixelout<=1'b1;
11603: pixelout<=1'b1;
11604: pixelout<=1'b1;
11605: pixelout<=1'b1;
11606: pixelout<=1'b1;
11607: pixelout<=1'b1;
11608: pixelout<=1'b1;
11609: pixelout<=1'b1;
11610: pixelout<=1'b1;
11611: pixelout<=1'b1;
11612: pixelout<=1'b1;
11613: pixelout<=1'b1;
11614: pixelout<=1'b1;
11615: pixelout<=1'b1;
11616: pixelout<=1'b1;
11617: pixelout<=1'b1;
11618: pixelout<=1'b1;
11619: pixelout<=1'b1;
11620: pixelout<=1'b1;
11621: pixelout<=1'b1;
11622: pixelout<=1'b1;
11623: pixelout<=1'b1;
11624: pixelout<=1'b1;
11625: pixelout<=1'b1;
11626: pixelout<=1'b1;
11627: pixelout<=1'b1;
11628: pixelout<=1'b1;
11629: pixelout<=1'b1;
11630: pixelout<=1'b1;
11631: pixelout<=1'b1;
11632: pixelout<=1'b1;
11633: pixelout<=1'b1;
11634: pixelout<=1'b1;
11635: pixelout<=1'b1;
11636: pixelout<=1'b1;
11637: pixelout<=1'b1;
11638: pixelout<=1'b1;
11639: pixelout<=1'b1;
11640: pixelout<=1'b1;
11641: pixelout<=1'b1;
11642: pixelout<=1'b1;
11643: pixelout<=1'b1;
11644: pixelout<=1'b1;
11645: pixelout<=1'b1;
11646: pixelout<=1'b1;
11647: pixelout<=1'b1;
11648: pixelout<=1'b1;
11649: pixelout<=1'b1;
11650: pixelout<=1'b1;
11651: pixelout<=1'b1;
11652: pixelout<=1'b1;
11653: pixelout<=1'b1;
11654: pixelout<=1'b1;
11655: pixelout<=1'b1;
11656: pixelout<=1'b1;
11657: pixelout<=1'b1;
11658: pixelout<=1'b1;
11659: pixelout<=1'b1;
11660: pixelout<=1'b1;
11661: pixelout<=1'b1;
11662: pixelout<=1'b1;
11663: pixelout<=1'b1;
11664: pixelout<=1'b1;
11665: pixelout<=1'b1;
11666: pixelout<=1'b1;
11667: pixelout<=1'b1;
11668: pixelout<=1'b1;
11669: pixelout<=1'b1;
11670: pixelout<=1'b1;
11671: pixelout<=1'b1;
11672: pixelout<=1'b1;
11673: pixelout<=1'b1;
11674: pixelout<=1'b1;
11675: pixelout<=1'b1;
11676: pixelout<=1'b1;
11677: pixelout<=1'b1;
11678: pixelout<=1'b1;
11679: pixelout<=1'b1;
11680: pixelout<=1'b1;
11681: pixelout<=1'b1;
11682: pixelout<=1'b1;
11683: pixelout<=1'b1;
11684: pixelout<=1'b1;
11685: pixelout<=1'b1;
11686: pixelout<=1'b1;
11687: pixelout<=1'b1;
11688: pixelout<=1'b1;
11689: pixelout<=1'b1;
11690: pixelout<=1'b1;
11691: pixelout<=1'b1;
11692: pixelout<=1'b1;
11693: pixelout<=1'b1;
11694: pixelout<=1'b1;
11695: pixelout<=1'b1;
11696: pixelout<=1'b1;
11697: pixelout<=1'b1;
11698: pixelout<=1'b1;
11699: pixelout<=1'b1;
11700: pixelout<=1'b1;
11701: pixelout<=1'b1;
11702: pixelout<=1'b1;
11703: pixelout<=1'b1;
11704: pixelout<=1'b1;
11705: pixelout<=1'b1;
11706: pixelout<=1'b1;
11707: pixelout<=1'b1;
11708: pixelout<=1'b1;
11709: pixelout<=1'b1;
11710: pixelout<=1'b1;
11711: pixelout<=1'b1;
11712: pixelout<=1'b1;
11713: pixelout<=1'b1;
11714: pixelout<=1'b1;
11715: pixelout<=1'b1;
11716: pixelout<=1'b1;
11717: pixelout<=1'b1;
11718: pixelout<=1'b1;
11719: pixelout<=1'b1;
11720: pixelout<=1'b1;
11721: pixelout<=1'b1;
11722: pixelout<=1'b1;
11723: pixelout<=1'b1;
11724: pixelout<=1'b1;
11725: pixelout<=1'b1;
11726: pixelout<=1'b1;
11727: pixelout<=1'b1;
11728: pixelout<=1'b1;
11729: pixelout<=1'b1;
11730: pixelout<=1'b1;
11731: pixelout<=1'b1;
11732: pixelout<=1'b1;
11733: pixelout<=1'b1;
11734: pixelout<=1'b1;
11735: pixelout<=1'b1;
11736: pixelout<=1'b1;
11737: pixelout<=1'b1;
11738: pixelout<=1'b1;
11739: pixelout<=1'b1;
11740: pixelout<=1'b1;
11741: pixelout<=1'b1;
11742: pixelout<=1'b1;
11743: pixelout<=1'b1;
11744: pixelout<=1'b1;
11745: pixelout<=1'b1;
11746: pixelout<=1'b1;
11747: pixelout<=1'b1;
11748: pixelout<=1'b1;
11749: pixelout<=1'b1;
11750: pixelout<=1'b1;
11751: pixelout<=1'b1;
11752: pixelout<=1'b1;
11753: pixelout<=1'b1;
11754: pixelout<=1'b1;
11755: pixelout<=1'b1;
11756: pixelout<=1'b1;
11757: pixelout<=1'b1;
11758: pixelout<=1'b1;
11759: pixelout<=1'b1;
11760: pixelout<=1'b1;
11761: pixelout<=1'b1;
11762: pixelout<=1'b1;
11763: pixelout<=1'b1;
11764: pixelout<=1'b1;
11765: pixelout<=1'b1;
11766: pixelout<=1'b1;
11767: pixelout<=1'b1;
11768: pixelout<=1'b1;
11769: pixelout<=1'b1;
11770: pixelout<=1'b1;
11771: pixelout<=1'b1;
11772: pixelout<=1'b1;
11773: pixelout<=1'b1;
11774: pixelout<=1'b1;
11775: pixelout<=1'b1;
11776: pixelout<=1'b1;
11777: pixelout<=1'b1;
11778: pixelout<=1'b1;
11779: pixelout<=1'b1;
11780: pixelout<=1'b1;
11781: pixelout<=1'b1;
11782: pixelout<=1'b1;
11783: pixelout<=1'b1;
11784: pixelout<=1'b1;
11785: pixelout<=1'b1;
11786: pixelout<=1'b1;
11787: pixelout<=1'b1;
11788: pixelout<=1'b1;
11789: pixelout<=1'b1;
11790: pixelout<=1'b1;
11791: pixelout<=1'b1;
11792: pixelout<=1'b1;
11793: pixelout<=1'b1;
11794: pixelout<=1'b1;
11795: pixelout<=1'b1;
11796: pixelout<=1'b1;
11797: pixelout<=1'b1;
11798: pixelout<=1'b1;
11799: pixelout<=1'b1;
11800: pixelout<=1'b1;
11801: pixelout<=1'b1;
11802: pixelout<=1'b1;
11803: pixelout<=1'b1;
11804: pixelout<=1'b1;
11805: pixelout<=1'b1;
11806: pixelout<=1'b1;
11807: pixelout<=1'b1;
11808: pixelout<=1'b1;
11809: pixelout<=1'b1;
11810: pixelout<=1'b1;
11811: pixelout<=1'b1;
11812: pixelout<=1'b1;
11813: pixelout<=1'b1;
11814: pixelout<=1'b1;
11815: pixelout<=1'b1;
11816: pixelout<=1'b1;
11817: pixelout<=1'b1;
11818: pixelout<=1'b1;
11819: pixelout<=1'b1;
11820: pixelout<=1'b1;
11821: pixelout<=1'b1;
11822: pixelout<=1'b1;
11823: pixelout<=1'b1;
11824: pixelout<=1'b1;
11825: pixelout<=1'b1;
11826: pixelout<=1'b1;
11827: pixelout<=1'b1;
11828: pixelout<=1'b1;
11829: pixelout<=1'b1;
11830: pixelout<=1'b1;
11831: pixelout<=1'b1;
11832: pixelout<=1'b1;
11833: pixelout<=1'b1;
11834: pixelout<=1'b1;
11835: pixelout<=1'b1;
11836: pixelout<=1'b1;
11837: pixelout<=1'b1;
11838: pixelout<=1'b1;
11839: pixelout<=1'b1;
11840: pixelout<=1'b1;
11841: pixelout<=1'b1;
11842: pixelout<=1'b1;
11843: pixelout<=1'b1;
11844: pixelout<=1'b1;
11845: pixelout<=1'b1;
11846: pixelout<=1'b1;
11847: pixelout<=1'b1;
11848: pixelout<=1'b1;
11849: pixelout<=1'b1;
11850: pixelout<=1'b1;
11851: pixelout<=1'b1;
11852: pixelout<=1'b1;
11853: pixelout<=1'b1;
11854: pixelout<=1'b1;
11855: pixelout<=1'b1;
11856: pixelout<=1'b1;
11857: pixelout<=1'b1;
11858: pixelout<=1'b1;
11859: pixelout<=1'b1;
11860: pixelout<=1'b1;
11861: pixelout<=1'b1;
11862: pixelout<=1'b1;
11863: pixelout<=1'b1;
11864: pixelout<=1'b1;
11865: pixelout<=1'b1;
11866: pixelout<=1'b1;
11867: pixelout<=1'b1;
11868: pixelout<=1'b1;
11869: pixelout<=1'b1;
11870: pixelout<=1'b1;
11871: pixelout<=1'b1;
11872: pixelout<=1'b1;
11873: pixelout<=1'b1;
11874: pixelout<=1'b1;
11875: pixelout<=1'b1;
11876: pixelout<=1'b1;
11877: pixelout<=1'b1;
11878: pixelout<=1'b1;
11879: pixelout<=1'b1;
11880: pixelout<=1'b1;
11881: pixelout<=1'b1;
11882: pixelout<=1'b1;
11883: pixelout<=1'b1;
11884: pixelout<=1'b1;
11885: pixelout<=1'b1;
11886: pixelout<=1'b1;
11887: pixelout<=1'b1;
11888: pixelout<=1'b1;
11889: pixelout<=1'b1;
11890: pixelout<=1'b1;
11891: pixelout<=1'b1;
11892: pixelout<=1'b1;
11893: pixelout<=1'b1;
11894: pixelout<=1'b1;
11895: pixelout<=1'b1;
11896: pixelout<=1'b1;
11897: pixelout<=1'b1;
11898: pixelout<=1'b1;
11899: pixelout<=1'b1;
11900: pixelout<=1'b1;
11901: pixelout<=1'b1;
11902: pixelout<=1'b1;
11903: pixelout<=1'b1;
11904: pixelout<=1'b1;
11905: pixelout<=1'b1;
11906: pixelout<=1'b1;
11907: pixelout<=1'b1;
11908: pixelout<=1'b1;
11909: pixelout<=1'b1;
11910: pixelout<=1'b1;
11911: pixelout<=1'b1;
11912: pixelout<=1'b1;
11913: pixelout<=1'b1;
11914: pixelout<=1'b1;
11915: pixelout<=1'b1;
11916: pixelout<=1'b1;
11917: pixelout<=1'b1;
11918: pixelout<=1'b1;
11919: pixelout<=1'b1;
11920: pixelout<=1'b1;
11921: pixelout<=1'b1;
11922: pixelout<=1'b1;
11923: pixelout<=1'b1;
11924: pixelout<=1'b1;
11925: pixelout<=1'b1;
11926: pixelout<=1'b1;
11927: pixelout<=1'b1;
11928: pixelout<=1'b1;
11929: pixelout<=1'b1;
11930: pixelout<=1'b1;
11931: pixelout<=1'b1;
11932: pixelout<=1'b1;
11933: pixelout<=1'b1;
11934: pixelout<=1'b1;
11935: pixelout<=1'b1;
11936: pixelout<=1'b1;
11937: pixelout<=1'b1;
11938: pixelout<=1'b1;
11939: pixelout<=1'b1;
11940: pixelout<=1'b1;
11941: pixelout<=1'b1;
11942: pixelout<=1'b1;
11943: pixelout<=1'b1;
11944: pixelout<=1'b1;
11945: pixelout<=1'b1;
11946: pixelout<=1'b1;
11947: pixelout<=1'b1;
11948: pixelout<=1'b1;
11949: pixelout<=1'b1;
11950: pixelout<=1'b1;
11951: pixelout<=1'b1;
11952: pixelout<=1'b1;
11953: pixelout<=1'b1;
11954: pixelout<=1'b1;
11955: pixelout<=1'b1;
11956: pixelout<=1'b1;
11957: pixelout<=1'b1;
11958: pixelout<=1'b1;
11959: pixelout<=1'b1;
11960: pixelout<=1'b1;
11961: pixelout<=1'b1;
11962: pixelout<=1'b1;
11963: pixelout<=1'b1;
11964: pixelout<=1'b1;
11965: pixelout<=1'b1;
11966: pixelout<=1'b1;
11967: pixelout<=1'b1;
11968: pixelout<=1'b1;
11969: pixelout<=1'b1;
11970: pixelout<=1'b1;
11971: pixelout<=1'b1;
11972: pixelout<=1'b1;
11973: pixelout<=1'b1;
11974: pixelout<=1'b1;
11975: pixelout<=1'b1;
11976: pixelout<=1'b1;
11977: pixelout<=1'b1;
11978: pixelout<=1'b1;
11979: pixelout<=1'b1;
11980: pixelout<=1'b1;
11981: pixelout<=1'b1;
11982: pixelout<=1'b1;
11983: pixelout<=1'b1;
11984: pixelout<=1'b1;
11985: pixelout<=1'b1;
11986: pixelout<=1'b1;
11987: pixelout<=1'b1;
11988: pixelout<=1'b1;
11989: pixelout<=1'b1;
11990: pixelout<=1'b1;
11991: pixelout<=1'b1;
11992: pixelout<=1'b1;
11993: pixelout<=1'b1;
11994: pixelout<=1'b1;
11995: pixelout<=1'b1;
11996: pixelout<=1'b1;
11997: pixelout<=1'b1;
11998: pixelout<=1'b1;
11999: pixelout<=1'b1;
12000: pixelout<=1'b1;
12001: pixelout<=1'b1;
12002: pixelout<=1'b1;
12003: pixelout<=1'b1;
12004: pixelout<=1'b1;
12005: pixelout<=1'b1;
12006: pixelout<=1'b1;
12007: pixelout<=1'b1;
12008: pixelout<=1'b1;
12009: pixelout<=1'b1;
12010: pixelout<=1'b1;
12011: pixelout<=1'b1;
12012: pixelout<=1'b1;
12013: pixelout<=1'b1;
12014: pixelout<=1'b1;
12015: pixelout<=1'b1;
12016: pixelout<=1'b1;
12017: pixelout<=1'b1;
12018: pixelout<=1'b1;
12019: pixelout<=1'b1;
12020: pixelout<=1'b1;
12021: pixelout<=1'b1;
12022: pixelout<=1'b1;
12023: pixelout<=1'b1;
12024: pixelout<=1'b1;
12025: pixelout<=1'b1;
12026: pixelout<=1'b1;
12027: pixelout<=1'b1;
12028: pixelout<=1'b1;
12029: pixelout<=1'b1;
12030: pixelout<=1'b1;
12031: pixelout<=1'b1;
12032: pixelout<=1'b1;
12033: pixelout<=1'b1;
12034: pixelout<=1'b1;
12035: pixelout<=1'b1;
12036: pixelout<=1'b1;
12037: pixelout<=1'b1;
12038: pixelout<=1'b1;
12039: pixelout<=1'b1;
12040: pixelout<=1'b1;
12041: pixelout<=1'b1;
12042: pixelout<=1'b1;
12043: pixelout<=1'b1;
12044: pixelout<=1'b1;
12045: pixelout<=1'b1;
12046: pixelout<=1'b1;
12047: pixelout<=1'b1;
12048: pixelout<=1'b1;
12049: pixelout<=1'b1;
12050: pixelout<=1'b1;
12051: pixelout<=1'b1;
12052: pixelout<=1'b1;
12053: pixelout<=1'b1;
12054: pixelout<=1'b1;
12055: pixelout<=1'b1;
12056: pixelout<=1'b1;
12057: pixelout<=1'b1;
12058: pixelout<=1'b1;
12059: pixelout<=1'b1;
12060: pixelout<=1'b1;
12061: pixelout<=1'b1;
12062: pixelout<=1'b1;
12063: pixelout<=1'b1;
12064: pixelout<=1'b1;
12065: pixelout<=1'b1;
12066: pixelout<=1'b1;
12067: pixelout<=1'b1;
12068: pixelout<=1'b1;
12069: pixelout<=1'b1;
12070: pixelout<=1'b1;
12071: pixelout<=1'b1;
12072: pixelout<=1'b1;
12073: pixelout<=1'b1;
12074: pixelout<=1'b1;
12075: pixelout<=1'b1;
12076: pixelout<=1'b1;
12077: pixelout<=1'b1;
12078: pixelout<=1'b1;
12079: pixelout<=1'b1;
12080: pixelout<=1'b1;
12081: pixelout<=1'b1;
12082: pixelout<=1'b1;
12083: pixelout<=1'b1;
12084: pixelout<=1'b1;
12085: pixelout<=1'b1;
12086: pixelout<=1'b1;
12087: pixelout<=1'b1;
12088: pixelout<=1'b1;
12089: pixelout<=1'b1;
12090: pixelout<=1'b1;
12091: pixelout<=1'b1;
12092: pixelout<=1'b1;
12093: pixelout<=1'b1;
12094: pixelout<=1'b1;
12095: pixelout<=1'b1;
12096: pixelout<=1'b1;
12097: pixelout<=1'b1;
12098: pixelout<=1'b1;
12099: pixelout<=1'b1;
12100: pixelout<=1'b1;
12101: pixelout<=1'b1;
12102: pixelout<=1'b1;
12103: pixelout<=1'b1;
12104: pixelout<=1'b1;
12105: pixelout<=1'b1;
12106: pixelout<=1'b1;
12107: pixelout<=1'b1;
12108: pixelout<=1'b1;
12109: pixelout<=1'b1;
12110: pixelout<=1'b1;
12111: pixelout<=1'b1;
12112: pixelout<=1'b1;
12113: pixelout<=1'b1;
12114: pixelout<=1'b1;
12115: pixelout<=1'b1;
12116: pixelout<=1'b1;
12117: pixelout<=1'b1;
12118: pixelout<=1'b1;
12119: pixelout<=1'b1;
12120: pixelout<=1'b1;
12121: pixelout<=1'b1;
12122: pixelout<=1'b1;
12123: pixelout<=1'b1;
12124: pixelout<=1'b1;
12125: pixelout<=1'b1;
12126: pixelout<=1'b1;
12127: pixelout<=1'b1;
12128: pixelout<=1'b1;
12129: pixelout<=1'b1;
12130: pixelout<=1'b1;
12131: pixelout<=1'b1;
12132: pixelout<=1'b1;
12133: pixelout<=1'b1;
12134: pixelout<=1'b1;
12135: pixelout<=1'b1;
12136: pixelout<=1'b1;
12137: pixelout<=1'b1;
12138: pixelout<=1'b1;
12139: pixelout<=1'b1;
12140: pixelout<=1'b1;
12141: pixelout<=1'b1;
12142: pixelout<=1'b1;
12143: pixelout<=1'b1;
12144: pixelout<=1'b1;
12145: pixelout<=1'b1;
12146: pixelout<=1'b1;
12147: pixelout<=1'b1;
12148: pixelout<=1'b1;
12149: pixelout<=1'b1;
12150: pixelout<=1'b1;
12151: pixelout<=1'b1;
12152: pixelout<=1'b1;
12153: pixelout<=1'b1;
12154: pixelout<=1'b1;
12155: pixelout<=1'b1;
12156: pixelout<=1'b1;
12157: pixelout<=1'b1;
12158: pixelout<=1'b1;
12159: pixelout<=1'b1;
12160: pixelout<=1'b1;
12161: pixelout<=1'b1;
12162: pixelout<=1'b1;
12163: pixelout<=1'b1;
12164: pixelout<=1'b1;
12165: pixelout<=1'b1;
12166: pixelout<=1'b1;
12167: pixelout<=1'b1;
12168: pixelout<=1'b1;
12169: pixelout<=1'b1;
12170: pixelout<=1'b1;
12171: pixelout<=1'b1;
12172: pixelout<=1'b1;
12173: pixelout<=1'b1;
12174: pixelout<=1'b1;
12175: pixelout<=1'b1;
12176: pixelout<=1'b1;
12177: pixelout<=1'b1;
12178: pixelout<=1'b1;
12179: pixelout<=1'b1;
12180: pixelout<=1'b1;
12181: pixelout<=1'b1;
12182: pixelout<=1'b1;
12183: pixelout<=1'b1;
12184: pixelout<=1'b1;
12185: pixelout<=1'b1;
12186: pixelout<=1'b1;
12187: pixelout<=1'b1;
12188: pixelout<=1'b1;
12189: pixelout<=1'b1;
12190: pixelout<=1'b1;
12191: pixelout<=1'b1;
12192: pixelout<=1'b1;
12193: pixelout<=1'b1;
12194: pixelout<=1'b1;
12195: pixelout<=1'b1;
12196: pixelout<=1'b1;
12197: pixelout<=1'b1;
12198: pixelout<=1'b1;
12199: pixelout<=1'b1;
12200: pixelout<=1'b1;
12201: pixelout<=1'b1;
12202: pixelout<=1'b1;
12203: pixelout<=1'b1;
12204: pixelout<=1'b1;
12205: pixelout<=1'b1;
12206: pixelout<=1'b1;
12207: pixelout<=1'b1;
12208: pixelout<=1'b1;
12209: pixelout<=1'b1;
12210: pixelout<=1'b1;
12211: pixelout<=1'b1;
12212: pixelout<=1'b1;
12213: pixelout<=1'b1;
12214: pixelout<=1'b1;
12215: pixelout<=1'b1;
12216: pixelout<=1'b1;
12217: pixelout<=1'b1;
12218: pixelout<=1'b1;
12219: pixelout<=1'b1;
12220: pixelout<=1'b1;
12221: pixelout<=1'b1;
12222: pixelout<=1'b1;
12223: pixelout<=1'b1;
12224: pixelout<=1'b1;
12225: pixelout<=1'b1;
12226: pixelout<=1'b1;
12227: pixelout<=1'b1;
12228: pixelout<=1'b1;
12229: pixelout<=1'b1;
12230: pixelout<=1'b1;
12231: pixelout<=1'b1;
12232: pixelout<=1'b1;
12233: pixelout<=1'b1;
12234: pixelout<=1'b1;
12235: pixelout<=1'b1;
12236: pixelout<=1'b1;
12237: pixelout<=1'b1;
12238: pixelout<=1'b1;
12239: pixelout<=1'b1;
12240: pixelout<=1'b1;
12241: pixelout<=1'b1;
12242: pixelout<=1'b1;
12243: pixelout<=1'b1;
12244: pixelout<=1'b1;
12245: pixelout<=1'b1;
12246: pixelout<=1'b1;
12247: pixelout<=1'b1;
12248: pixelout<=1'b1;
12249: pixelout<=1'b1;
12250: pixelout<=1'b1;
12251: pixelout<=1'b1;
12252: pixelout<=1'b1;
12253: pixelout<=1'b1;
12254: pixelout<=1'b1;
12255: pixelout<=1'b1;
12256: pixelout<=1'b1;
12257: pixelout<=1'b1;
12258: pixelout<=1'b1;
12259: pixelout<=1'b1;
12260: pixelout<=1'b1;
12261: pixelout<=1'b1;
12262: pixelout<=1'b1;
12263: pixelout<=1'b1;
12264: pixelout<=1'b1;
12265: pixelout<=1'b1;
12266: pixelout<=1'b1;
12267: pixelout<=1'b1;
12268: pixelout<=1'b1;
12269: pixelout<=1'b1;
12270: pixelout<=1'b1;
12271: pixelout<=1'b0;
12272: pixelout<=1'b0;
12273: pixelout<=1'b1;
12274: pixelout<=1'b1;
12275: pixelout<=1'b1;
12276: pixelout<=1'b1;
12277: pixelout<=1'b1;
12278: pixelout<=1'b1;
12279: pixelout<=1'b1;
12280: pixelout<=1'b1;
12281: pixelout<=1'b1;
12282: pixelout<=1'b1;
12283: pixelout<=1'b1;
12284: pixelout<=1'b1;
12285: pixelout<=1'b1;
12286: pixelout<=1'b1;
12287: pixelout<=1'b1;
12288: pixelout<=1'b1;
12289: pixelout<=1'b1;
12290: pixelout<=1'b1;
12291: pixelout<=1'b1;
12292: pixelout<=1'b1;
12293: pixelout<=1'b1;
12294: pixelout<=1'b1;
12295: pixelout<=1'b1;
12296: pixelout<=1'b1;
12297: pixelout<=1'b1;
12298: pixelout<=1'b1;
12299: pixelout<=1'b1;
12300: pixelout<=1'b1;
12301: pixelout<=1'b1;
12302: pixelout<=1'b1;
12303: pixelout<=1'b0;
12304: pixelout<=1'b1;
12305: pixelout<=1'b1;
12306: pixelout<=1'b1;
12307: pixelout<=1'b1;
12308: pixelout<=1'b1;
12309: pixelout<=1'b1;
12310: pixelout<=1'b1;
12311: pixelout<=1'b1;
12312: pixelout<=1'b1;
12313: pixelout<=1'b0;
12314: pixelout<=1'b1;
12315: pixelout<=1'b1;
12316: pixelout<=1'b1;
12317: pixelout<=1'b1;
12318: pixelout<=1'b1;
12319: pixelout<=1'b1;
12320: pixelout<=1'b1;
12321: pixelout<=1'b1;
12322: pixelout<=1'b1;
12323: pixelout<=1'b1;
12324: pixelout<=1'b1;
12325: pixelout<=1'b1;
12326: pixelout<=1'b1;
12327: pixelout<=1'b1;
12328: pixelout<=1'b1;
12329: pixelout<=1'b1;
12330: pixelout<=1'b1;
12331: pixelout<=1'b0;
12332: pixelout<=1'b1;
12333: pixelout<=1'b1;
12334: pixelout<=1'b1;
12335: pixelout<=1'b1;
12336: pixelout<=1'b1;
12337: pixelout<=1'b1;
12338: pixelout<=1'b1;
12339: pixelout<=1'b1;
12340: pixelout<=1'b1;
12341: pixelout<=1'b1;
12342: pixelout<=1'b1;
12343: pixelout<=1'b1;
12344: pixelout<=1'b1;
12345: pixelout<=1'b1;
12346: pixelout<=1'b1;
12347: pixelout<=1'b1;
12348: pixelout<=1'b1;
12349: pixelout<=1'b1;
12350: pixelout<=1'b1;
12351: pixelout<=1'b1;
12352: pixelout<=1'b1;
12353: pixelout<=1'b1;
12354: pixelout<=1'b1;
12355: pixelout<=1'b1;
12356: pixelout<=1'b1;
12357: pixelout<=1'b1;
12358: pixelout<=1'b1;
12359: pixelout<=1'b1;
12360: pixelout<=1'b1;
12361: pixelout<=1'b1;
12362: pixelout<=1'b1;
12363: pixelout<=1'b1;
12364: pixelout<=1'b1;
12365: pixelout<=1'b1;
12366: pixelout<=1'b1;
12367: pixelout<=1'b1;
12368: pixelout<=1'b1;
12369: pixelout<=1'b1;
12370: pixelout<=1'b1;
12371: pixelout<=1'b1;
12372: pixelout<=1'b1;
12373: pixelout<=1'b1;
12374: pixelout<=1'b1;
12375: pixelout<=1'b1;
12376: pixelout<=1'b1;
12377: pixelout<=1'b0;
12378: pixelout<=1'b0;
12379: pixelout<=1'b0;
12380: pixelout<=1'b0;
12381: pixelout<=1'b1;
12382: pixelout<=1'b1;
12383: pixelout<=1'b1;
12384: pixelout<=1'b0;
12385: pixelout<=1'b0;
12386: pixelout<=1'b0;
12387: pixelout<=1'b1;
12388: pixelout<=1'b1;
12389: pixelout<=1'b1;
12390: pixelout<=1'b1;
12391: pixelout<=1'b0;
12392: pixelout<=1'b0;
12393: pixelout<=1'b0;
12394: pixelout<=1'b0;
12395: pixelout<=1'b1;
12396: pixelout<=1'b1;
12397: pixelout<=1'b1;
12398: pixelout<=1'b1;
12399: pixelout<=1'b1;
12400: pixelout<=1'b1;
12401: pixelout<=1'b1;
12402: pixelout<=1'b1;
12403: pixelout<=1'b1;
12404: pixelout<=1'b1;
12405: pixelout<=1'b1;
12406: pixelout<=1'b1;
12407: pixelout<=1'b1;
12408: pixelout<=1'b1;
12409: pixelout<=1'b1;
12410: pixelout<=1'b1;
12411: pixelout<=1'b1;
12412: pixelout<=1'b1;
12413: pixelout<=1'b1;
12414: pixelout<=1'b1;
12415: pixelout<=1'b1;
12416: pixelout<=1'b1;
12417: pixelout<=1'b1;
12418: pixelout<=1'b1;
12419: pixelout<=1'b1;
12420: pixelout<=1'b1;
12421: pixelout<=1'b1;
12422: pixelout<=1'b1;
12423: pixelout<=1'b1;
12424: pixelout<=1'b1;
12425: pixelout<=1'b1;
12426: pixelout<=1'b1;
12427: pixelout<=1'b1;
12428: pixelout<=1'b1;
12429: pixelout<=1'b1;
12430: pixelout<=1'b1;
12431: pixelout<=1'b1;
12432: pixelout<=1'b1;
12433: pixelout<=1'b1;
12434: pixelout<=1'b1;
12435: pixelout<=1'b1;
12436: pixelout<=1'b1;
12437: pixelout<=1'b1;
12438: pixelout<=1'b1;
12439: pixelout<=1'b1;
12440: pixelout<=1'b1;
12441: pixelout<=1'b1;
12442: pixelout<=1'b1;
12443: pixelout<=1'b1;
12444: pixelout<=1'b1;
12445: pixelout<=1'b1;
12446: pixelout<=1'b1;
12447: pixelout<=1'b1;
12448: pixelout<=1'b1;
12449: pixelout<=1'b1;
12450: pixelout<=1'b1;
12451: pixelout<=1'b1;
12452: pixelout<=1'b1;
12453: pixelout<=1'b1;
12454: pixelout<=1'b1;
12455: pixelout<=1'b1;
12456: pixelout<=1'b1;
12457: pixelout<=1'b1;
12458: pixelout<=1'b1;
12459: pixelout<=1'b1;
12460: pixelout<=1'b1;
12461: pixelout<=1'b1;
12462: pixelout<=1'b1;
12463: pixelout<=1'b1;
12464: pixelout<=1'b1;
12465: pixelout<=1'b1;
12466: pixelout<=1'b1;
12467: pixelout<=1'b1;
12468: pixelout<=1'b1;
12469: pixelout<=1'b1;
12470: pixelout<=1'b1;
12471: pixelout<=1'b1;
12472: pixelout<=1'b1;
12473: pixelout<=1'b1;
12474: pixelout<=1'b1;
12475: pixelout<=1'b1;
12476: pixelout<=1'b1;
12477: pixelout<=1'b1;
12478: pixelout<=1'b1;
12479: pixelout<=1'b1;
12480: pixelout<=1'b1;
12481: pixelout<=1'b1;
12482: pixelout<=1'b1;
12483: pixelout<=1'b1;
12484: pixelout<=1'b1;
12485: pixelout<=1'b1;
12486: pixelout<=1'b1;
12487: pixelout<=1'b1;
12488: pixelout<=1'b1;
12489: pixelout<=1'b1;
12490: pixelout<=1'b1;
12491: pixelout<=1'b1;
12492: pixelout<=1'b1;
12493: pixelout<=1'b1;
12494: pixelout<=1'b1;
12495: pixelout<=1'b1;
12496: pixelout<=1'b1;
12497: pixelout<=1'b1;
12498: pixelout<=1'b1;
12499: pixelout<=1'b1;
12500: pixelout<=1'b1;
12501: pixelout<=1'b1;
12502: pixelout<=1'b1;
12503: pixelout<=1'b1;
12504: pixelout<=1'b1;
12505: pixelout<=1'b1;
12506: pixelout<=1'b1;
12507: pixelout<=1'b1;
12508: pixelout<=1'b1;
12509: pixelout<=1'b0;
12510: pixelout<=1'b1;
12511: pixelout<=1'b1;
12512: pixelout<=1'b1;
12513: pixelout<=1'b1;
12514: pixelout<=1'b1;
12515: pixelout<=1'b1;
12516: pixelout<=1'b1;
12517: pixelout<=1'b1;
12518: pixelout<=1'b1;
12519: pixelout<=1'b1;
12520: pixelout<=1'b1;
12521: pixelout<=1'b1;
12522: pixelout<=1'b1;
12523: pixelout<=1'b1;
12524: pixelout<=1'b1;
12525: pixelout<=1'b1;
12526: pixelout<=1'b1;
12527: pixelout<=1'b1;
12528: pixelout<=1'b1;
12529: pixelout<=1'b1;
12530: pixelout<=1'b1;
12531: pixelout<=1'b1;
12532: pixelout<=1'b1;
12533: pixelout<=1'b1;
12534: pixelout<=1'b1;
12535: pixelout<=1'b1;
12536: pixelout<=1'b1;
12537: pixelout<=1'b1;
12538: pixelout<=1'b1;
12539: pixelout<=1'b1;
12540: pixelout<=1'b1;
12541: pixelout<=1'b1;
12542: pixelout<=1'b1;
12543: pixelout<=1'b1;
12544: pixelout<=1'b1;
12545: pixelout<=1'b1;
12546: pixelout<=1'b1;
12547: pixelout<=1'b1;
12548: pixelout<=1'b1;
12549: pixelout<=1'b0;
12550: pixelout<=1'b1;
12551: pixelout<=1'b1;
12552: pixelout<=1'b1;
12553: pixelout<=1'b0;
12554: pixelout<=1'b1;
12555: pixelout<=1'b1;
12556: pixelout<=1'b1;
12557: pixelout<=1'b1;
12558: pixelout<=1'b1;
12559: pixelout<=1'b1;
12560: pixelout<=1'b1;
12561: pixelout<=1'b1;
12562: pixelout<=1'b1;
12563: pixelout<=1'b1;
12564: pixelout<=1'b1;
12565: pixelout<=1'b1;
12566: pixelout<=1'b1;
12567: pixelout<=1'b1;
12568: pixelout<=1'b1;
12569: pixelout<=1'b1;
12570: pixelout<=1'b1;
12571: pixelout<=1'b0;
12572: pixelout<=1'b1;
12573: pixelout<=1'b1;
12574: pixelout<=1'b1;
12575: pixelout<=1'b1;
12576: pixelout<=1'b1;
12577: pixelout<=1'b1;
12578: pixelout<=1'b1;
12579: pixelout<=1'b1;
12580: pixelout<=1'b1;
12581: pixelout<=1'b1;
12582: pixelout<=1'b1;
12583: pixelout<=1'b1;
12584: pixelout<=1'b0;
12585: pixelout<=1'b1;
12586: pixelout<=1'b1;
12587: pixelout<=1'b1;
12588: pixelout<=1'b1;
12589: pixelout<=1'b1;
12590: pixelout<=1'b1;
12591: pixelout<=1'b1;
12592: pixelout<=1'b1;
12593: pixelout<=1'b1;
12594: pixelout<=1'b1;
12595: pixelout<=1'b1;
12596: pixelout<=1'b1;
12597: pixelout<=1'b1;
12598: pixelout<=1'b1;
12599: pixelout<=1'b1;
12600: pixelout<=1'b1;
12601: pixelout<=1'b1;
12602: pixelout<=1'b1;
12603: pixelout<=1'b1;
12604: pixelout<=1'b1;
12605: pixelout<=1'b1;
12606: pixelout<=1'b1;
12607: pixelout<=1'b1;
12608: pixelout<=1'b1;
12609: pixelout<=1'b1;
12610: pixelout<=1'b1;
12611: pixelout<=1'b1;
12612: pixelout<=1'b1;
12613: pixelout<=1'b1;
12614: pixelout<=1'b1;
12615: pixelout<=1'b1;
12616: pixelout<=1'b1;
12617: pixelout<=1'b1;
12618: pixelout<=1'b1;
12619: pixelout<=1'b0;
12620: pixelout<=1'b1;
12621: pixelout<=1'b1;
12622: pixelout<=1'b1;
12623: pixelout<=1'b0;
12624: pixelout<=1'b1;
12625: pixelout<=1'b1;
12626: pixelout<=1'b1;
12627: pixelout<=1'b0;
12628: pixelout<=1'b1;
12629: pixelout<=1'b1;
12630: pixelout<=1'b1;
12631: pixelout<=1'b0;
12632: pixelout<=1'b1;
12633: pixelout<=1'b1;
12634: pixelout<=1'b1;
12635: pixelout<=1'b0;
12636: pixelout<=1'b1;
12637: pixelout<=1'b1;
12638: pixelout<=1'b1;
12639: pixelout<=1'b1;
12640: pixelout<=1'b1;
12641: pixelout<=1'b1;
12642: pixelout<=1'b1;
12643: pixelout<=1'b1;
12644: pixelout<=1'b1;
12645: pixelout<=1'b1;
12646: pixelout<=1'b1;
12647: pixelout<=1'b1;
12648: pixelout<=1'b1;
12649: pixelout<=1'b1;
12650: pixelout<=1'b1;
12651: pixelout<=1'b1;
12652: pixelout<=1'b1;
12653: pixelout<=1'b1;
12654: pixelout<=1'b1;
12655: pixelout<=1'b1;
12656: pixelout<=1'b1;
12657: pixelout<=1'b1;
12658: pixelout<=1'b1;
12659: pixelout<=1'b1;
12660: pixelout<=1'b1;
12661: pixelout<=1'b1;
12662: pixelout<=1'b1;
12663: pixelout<=1'b1;
12664: pixelout<=1'b1;
12665: pixelout<=1'b1;
12666: pixelout<=1'b1;
12667: pixelout<=1'b1;
12668: pixelout<=1'b1;
12669: pixelout<=1'b1;
12670: pixelout<=1'b1;
12671: pixelout<=1'b1;
12672: pixelout<=1'b1;
12673: pixelout<=1'b1;
12674: pixelout<=1'b1;
12675: pixelout<=1'b1;
12676: pixelout<=1'b1;
12677: pixelout<=1'b1;
12678: pixelout<=1'b1;
12679: pixelout<=1'b1;
12680: pixelout<=1'b1;
12681: pixelout<=1'b1;
12682: pixelout<=1'b1;
12683: pixelout<=1'b1;
12684: pixelout<=1'b1;
12685: pixelout<=1'b1;
12686: pixelout<=1'b1;
12687: pixelout<=1'b1;
12688: pixelout<=1'b1;
12689: pixelout<=1'b1;
12690: pixelout<=1'b1;
12691: pixelout<=1'b1;
12692: pixelout<=1'b1;
12693: pixelout<=1'b1;
12694: pixelout<=1'b1;
12695: pixelout<=1'b1;
12696: pixelout<=1'b1;
12697: pixelout<=1'b1;
12698: pixelout<=1'b1;
12699: pixelout<=1'b1;
12700: pixelout<=1'b1;
12701: pixelout<=1'b1;
12702: pixelout<=1'b1;
12703: pixelout<=1'b1;
12704: pixelout<=1'b1;
12705: pixelout<=1'b1;
12706: pixelout<=1'b1;
12707: pixelout<=1'b1;
12708: pixelout<=1'b1;
12709: pixelout<=1'b1;
12710: pixelout<=1'b1;
12711: pixelout<=1'b1;
12712: pixelout<=1'b1;
12713: pixelout<=1'b1;
12714: pixelout<=1'b1;
12715: pixelout<=1'b1;
12716: pixelout<=1'b1;
12717: pixelout<=1'b1;
12718: pixelout<=1'b1;
12719: pixelout<=1'b1;
12720: pixelout<=1'b1;
12721: pixelout<=1'b1;
12722: pixelout<=1'b1;
12723: pixelout<=1'b1;
12724: pixelout<=1'b1;
12725: pixelout<=1'b1;
12726: pixelout<=1'b1;
12727: pixelout<=1'b1;
12728: pixelout<=1'b1;
12729: pixelout<=1'b1;
12730: pixelout<=1'b1;
12731: pixelout<=1'b1;
12732: pixelout<=1'b1;
12733: pixelout<=1'b1;
12734: pixelout<=1'b1;
12735: pixelout<=1'b1;
12736: pixelout<=1'b1;
12737: pixelout<=1'b1;
12738: pixelout<=1'b1;
12739: pixelout<=1'b1;
12740: pixelout<=1'b1;
12741: pixelout<=1'b1;
12742: pixelout<=1'b1;
12743: pixelout<=1'b1;
12744: pixelout<=1'b1;
12745: pixelout<=1'b1;
12746: pixelout<=1'b1;
12747: pixelout<=1'b1;
12748: pixelout<=1'b1;
12749: pixelout<=1'b1;
12750: pixelout<=1'b1;
12751: pixelout<=1'b1;
12752: pixelout<=1'b1;
12753: pixelout<=1'b1;
12754: pixelout<=1'b1;
12755: pixelout<=1'b1;
12756: pixelout<=1'b1;
12757: pixelout<=1'b1;
12758: pixelout<=1'b1;
12759: pixelout<=1'b1;
12760: pixelout<=1'b1;
12761: pixelout<=1'b1;
12762: pixelout<=1'b1;
12763: pixelout<=1'b1;
12764: pixelout<=1'b1;
12765: pixelout<=1'b1;
12766: pixelout<=1'b1;
12767: pixelout<=1'b1;
12768: pixelout<=1'b1;
12769: pixelout<=1'b1;
12770: pixelout<=1'b1;
12771: pixelout<=1'b1;
12772: pixelout<=1'b1;
12773: pixelout<=1'b1;
12774: pixelout<=1'b1;
12775: pixelout<=1'b1;
12776: pixelout<=1'b1;
12777: pixelout<=1'b1;
12778: pixelout<=1'b1;
12779: pixelout<=1'b1;
12780: pixelout<=1'b1;
12781: pixelout<=1'b1;
12782: pixelout<=1'b1;
12783: pixelout<=1'b1;
12784: pixelout<=1'b1;
12785: pixelout<=1'b1;
12786: pixelout<=1'b1;
12787: pixelout<=1'b1;
12788: pixelout<=1'b1;
12789: pixelout<=1'b0;
12790: pixelout<=1'b1;
12791: pixelout<=1'b1;
12792: pixelout<=1'b1;
12793: pixelout<=1'b0;
12794: pixelout<=1'b1;
12795: pixelout<=1'b1;
12796: pixelout<=1'b1;
12797: pixelout<=1'b1;
12798: pixelout<=1'b1;
12799: pixelout<=1'b1;
12800: pixelout<=1'b1;
12801: pixelout<=1'b1;
12802: pixelout<=1'b1;
12803: pixelout<=1'b1;
12804: pixelout<=1'b1;
12805: pixelout<=1'b1;
12806: pixelout<=1'b1;
12807: pixelout<=1'b1;
12808: pixelout<=1'b1;
12809: pixelout<=1'b1;
12810: pixelout<=1'b1;
12811: pixelout<=1'b0;
12812: pixelout<=1'b1;
12813: pixelout<=1'b1;
12814: pixelout<=1'b1;
12815: pixelout<=1'b1;
12816: pixelout<=1'b1;
12817: pixelout<=1'b1;
12818: pixelout<=1'b1;
12819: pixelout<=1'b1;
12820: pixelout<=1'b1;
12821: pixelout<=1'b1;
12822: pixelout<=1'b1;
12823: pixelout<=1'b1;
12824: pixelout<=1'b0;
12825: pixelout<=1'b1;
12826: pixelout<=1'b1;
12827: pixelout<=1'b1;
12828: pixelout<=1'b1;
12829: pixelout<=1'b1;
12830: pixelout<=1'b1;
12831: pixelout<=1'b1;
12832: pixelout<=1'b1;
12833: pixelout<=1'b1;
12834: pixelout<=1'b1;
12835: pixelout<=1'b1;
12836: pixelout<=1'b1;
12837: pixelout<=1'b1;
12838: pixelout<=1'b1;
12839: pixelout<=1'b1;
12840: pixelout<=1'b1;
12841: pixelout<=1'b1;
12842: pixelout<=1'b1;
12843: pixelout<=1'b1;
12844: pixelout<=1'b1;
12845: pixelout<=1'b1;
12846: pixelout<=1'b1;
12847: pixelout<=1'b1;
12848: pixelout<=1'b1;
12849: pixelout<=1'b1;
12850: pixelout<=1'b1;
12851: pixelout<=1'b1;
12852: pixelout<=1'b1;
12853: pixelout<=1'b1;
12854: pixelout<=1'b1;
12855: pixelout<=1'b1;
12856: pixelout<=1'b1;
12857: pixelout<=1'b1;
12858: pixelout<=1'b1;
12859: pixelout<=1'b0;
12860: pixelout<=1'b1;
12861: pixelout<=1'b1;
12862: pixelout<=1'b1;
12863: pixelout<=1'b0;
12864: pixelout<=1'b1;
12865: pixelout<=1'b1;
12866: pixelout<=1'b1;
12867: pixelout<=1'b0;
12868: pixelout<=1'b1;
12869: pixelout<=1'b1;
12870: pixelout<=1'b1;
12871: pixelout<=1'b0;
12872: pixelout<=1'b1;
12873: pixelout<=1'b1;
12874: pixelout<=1'b1;
12875: pixelout<=1'b0;
12876: pixelout<=1'b1;
12877: pixelout<=1'b1;
12878: pixelout<=1'b1;
12879: pixelout<=1'b1;
12880: pixelout<=1'b1;
12881: pixelout<=1'b1;
12882: pixelout<=1'b1;
12883: pixelout<=1'b1;
12884: pixelout<=1'b1;
12885: pixelout<=1'b1;
12886: pixelout<=1'b1;
12887: pixelout<=1'b1;
12888: pixelout<=1'b1;
12889: pixelout<=1'b1;
12890: pixelout<=1'b1;
12891: pixelout<=1'b1;
12892: pixelout<=1'b1;
12893: pixelout<=1'b1;
12894: pixelout<=1'b1;
12895: pixelout<=1'b1;
12896: pixelout<=1'b1;
12897: pixelout<=1'b1;
12898: pixelout<=1'b1;
12899: pixelout<=1'b1;
12900: pixelout<=1'b1;
12901: pixelout<=1'b1;
12902: pixelout<=1'b1;
12903: pixelout<=1'b1;
12904: pixelout<=1'b1;
12905: pixelout<=1'b1;
12906: pixelout<=1'b1;
12907: pixelout<=1'b1;
12908: pixelout<=1'b1;
12909: pixelout<=1'b1;
12910: pixelout<=1'b1;
12911: pixelout<=1'b1;
12912: pixelout<=1'b1;
12913: pixelout<=1'b1;
12914: pixelout<=1'b1;
12915: pixelout<=1'b1;
12916: pixelout<=1'b1;
12917: pixelout<=1'b1;
12918: pixelout<=1'b1;
12919: pixelout<=1'b1;
12920: pixelout<=1'b1;
12921: pixelout<=1'b1;
12922: pixelout<=1'b1;
12923: pixelout<=1'b1;
12924: pixelout<=1'b1;
12925: pixelout<=1'b1;
12926: pixelout<=1'b1;
12927: pixelout<=1'b1;
12928: pixelout<=1'b1;
12929: pixelout<=1'b1;
12930: pixelout<=1'b1;
12931: pixelout<=1'b1;
12932: pixelout<=1'b1;
12933: pixelout<=1'b1;
12934: pixelout<=1'b1;
12935: pixelout<=1'b1;
12936: pixelout<=1'b1;
12937: pixelout<=1'b1;
12938: pixelout<=1'b1;
12939: pixelout<=1'b1;
12940: pixelout<=1'b1;
12941: pixelout<=1'b1;
12942: pixelout<=1'b1;
12943: pixelout<=1'b1;
12944: pixelout<=1'b1;
12945: pixelout<=1'b1;
12946: pixelout<=1'b1;
12947: pixelout<=1'b1;
12948: pixelout<=1'b1;
12949: pixelout<=1'b1;
12950: pixelout<=1'b1;
12951: pixelout<=1'b1;
12952: pixelout<=1'b1;
12953: pixelout<=1'b1;
12954: pixelout<=1'b1;
12955: pixelout<=1'b1;
12956: pixelout<=1'b1;
12957: pixelout<=1'b1;
12958: pixelout<=1'b1;
12959: pixelout<=1'b1;
12960: pixelout<=1'b1;
12961: pixelout<=1'b1;
12962: pixelout<=1'b1;
12963: pixelout<=1'b1;
12964: pixelout<=1'b1;
12965: pixelout<=1'b1;
12966: pixelout<=1'b1;
12967: pixelout<=1'b1;
12968: pixelout<=1'b1;
12969: pixelout<=1'b1;
12970: pixelout<=1'b1;
12971: pixelout<=1'b1;
12972: pixelout<=1'b1;
12973: pixelout<=1'b1;
12974: pixelout<=1'b1;
12975: pixelout<=1'b1;
12976: pixelout<=1'b1;
12977: pixelout<=1'b1;
12978: pixelout<=1'b1;
12979: pixelout<=1'b1;
12980: pixelout<=1'b1;
12981: pixelout<=1'b1;
12982: pixelout<=1'b1;
12983: pixelout<=1'b1;
12984: pixelout<=1'b1;
12985: pixelout<=1'b1;
12986: pixelout<=1'b1;
12987: pixelout<=1'b1;
12988: pixelout<=1'b1;
12989: pixelout<=1'b1;
12990: pixelout<=1'b1;
12991: pixelout<=1'b0;
12992: pixelout<=1'b1;
12993: pixelout<=1'b1;
12994: pixelout<=1'b1;
12995: pixelout<=1'b1;
12996: pixelout<=1'b0;
12997: pixelout<=1'b0;
12998: pixelout<=1'b0;
12999: pixelout<=1'b1;
13000: pixelout<=1'b1;
13001: pixelout<=1'b1;
13002: pixelout<=1'b1;
13003: pixelout<=1'b0;
13004: pixelout<=1'b0;
13005: pixelout<=1'b0;
13006: pixelout<=1'b1;
13007: pixelout<=1'b1;
13008: pixelout<=1'b1;
13009: pixelout<=1'b0;
13010: pixelout<=1'b0;
13011: pixelout<=1'b0;
13012: pixelout<=1'b1;
13013: pixelout<=1'b1;
13014: pixelout<=1'b0;
13015: pixelout<=1'b1;
13016: pixelout<=1'b1;
13017: pixelout<=1'b1;
13018: pixelout<=1'b0;
13019: pixelout<=1'b0;
13020: pixelout<=1'b0;
13021: pixelout<=1'b1;
13022: pixelout<=1'b1;
13023: pixelout<=1'b1;
13024: pixelout<=1'b1;
13025: pixelout<=1'b1;
13026: pixelout<=1'b1;
13027: pixelout<=1'b1;
13028: pixelout<=1'b0;
13029: pixelout<=1'b0;
13030: pixelout<=1'b0;
13031: pixelout<=1'b0;
13032: pixelout<=1'b1;
13033: pixelout<=1'b0;
13034: pixelout<=1'b0;
13035: pixelout<=1'b0;
13036: pixelout<=1'b0;
13037: pixelout<=1'b1;
13038: pixelout<=1'b1;
13039: pixelout<=1'b1;
13040: pixelout<=1'b1;
13041: pixelout<=1'b0;
13042: pixelout<=1'b0;
13043: pixelout<=1'b0;
13044: pixelout<=1'b1;
13045: pixelout<=1'b1;
13046: pixelout<=1'b0;
13047: pixelout<=1'b0;
13048: pixelout<=1'b1;
13049: pixelout<=1'b1;
13050: pixelout<=1'b1;
13051: pixelout<=1'b0;
13052: pixelout<=1'b1;
13053: pixelout<=1'b1;
13054: pixelout<=1'b0;
13055: pixelout<=1'b1;
13056: pixelout<=1'b0;
13057: pixelout<=1'b0;
13058: pixelout<=1'b0;
13059: pixelout<=1'b0;
13060: pixelout<=1'b1;
13061: pixelout<=1'b1;
13062: pixelout<=1'b1;
13063: pixelout<=1'b1;
13064: pixelout<=1'b0;
13065: pixelout<=1'b0;
13066: pixelout<=1'b0;
13067: pixelout<=1'b1;
13068: pixelout<=1'b1;
13069: pixelout<=1'b1;
13070: pixelout<=1'b0;
13071: pixelout<=1'b0;
13072: pixelout<=1'b1;
13073: pixelout<=1'b1;
13074: pixelout<=1'b1;
13075: pixelout<=1'b1;
13076: pixelout<=1'b1;
13077: pixelout<=1'b1;
13078: pixelout<=1'b0;
13079: pixelout<=1'b0;
13080: pixelout<=1'b0;
13081: pixelout<=1'b1;
13082: pixelout<=1'b1;
13083: pixelout<=1'b0;
13084: pixelout<=1'b1;
13085: pixelout<=1'b1;
13086: pixelout<=1'b0;
13087: pixelout<=1'b1;
13088: pixelout<=1'b1;
13089: pixelout<=1'b0;
13090: pixelout<=1'b1;
13091: pixelout<=1'b1;
13092: pixelout<=1'b0;
13093: pixelout<=1'b1;
13094: pixelout<=1'b1;
13095: pixelout<=1'b1;
13096: pixelout<=1'b1;
13097: pixelout<=1'b1;
13098: pixelout<=1'b1;
13099: pixelout<=1'b0;
13100: pixelout<=1'b1;
13101: pixelout<=1'b1;
13102: pixelout<=1'b1;
13103: pixelout<=1'b0;
13104: pixelout<=1'b1;
13105: pixelout<=1'b1;
13106: pixelout<=1'b1;
13107: pixelout<=1'b0;
13108: pixelout<=1'b1;
13109: pixelout<=1'b1;
13110: pixelout<=1'b1;
13111: pixelout<=1'b0;
13112: pixelout<=1'b1;
13113: pixelout<=1'b1;
13114: pixelout<=1'b1;
13115: pixelout<=1'b0;
13116: pixelout<=1'b1;
13117: pixelout<=1'b1;
13118: pixelout<=1'b1;
13119: pixelout<=1'b0;
13120: pixelout<=1'b0;
13121: pixelout<=1'b1;
13122: pixelout<=1'b1;
13123: pixelout<=1'b1;
13124: pixelout<=1'b0;
13125: pixelout<=1'b0;
13126: pixelout<=1'b0;
13127: pixelout<=1'b1;
13128: pixelout<=1'b1;
13129: pixelout<=1'b1;
13130: pixelout<=1'b0;
13131: pixelout<=1'b1;
13132: pixelout<=1'b1;
13133: pixelout<=1'b0;
13134: pixelout<=1'b1;
13135: pixelout<=1'b1;
13136: pixelout<=1'b0;
13137: pixelout<=1'b0;
13138: pixelout<=1'b0;
13139: pixelout<=1'b1;
13140: pixelout<=1'b1;
13141: pixelout<=1'b1;
13142: pixelout<=1'b1;
13143: pixelout<=1'b1;
13144: pixelout<=1'b1;
13145: pixelout<=1'b1;
13146: pixelout<=1'b1;
13147: pixelout<=1'b1;
13148: pixelout<=1'b1;
13149: pixelout<=1'b1;
13150: pixelout<=1'b1;
13151: pixelout<=1'b0;
13152: pixelout<=1'b0;
13153: pixelout<=1'b1;
13154: pixelout<=1'b1;
13155: pixelout<=1'b1;
13156: pixelout<=1'b1;
13157: pixelout<=1'b0;
13158: pixelout<=1'b0;
13159: pixelout<=1'b0;
13160: pixelout<=1'b1;
13161: pixelout<=1'b1;
13162: pixelout<=1'b0;
13163: pixelout<=1'b0;
13164: pixelout<=1'b0;
13165: pixelout<=1'b1;
13166: pixelout<=1'b1;
13167: pixelout<=1'b1;
13168: pixelout<=1'b1;
13169: pixelout<=1'b1;
13170: pixelout<=1'b1;
13171: pixelout<=1'b1;
13172: pixelout<=1'b1;
13173: pixelout<=1'b1;
13174: pixelout<=1'b1;
13175: pixelout<=1'b1;
13176: pixelout<=1'b1;
13177: pixelout<=1'b1;
13178: pixelout<=1'b1;
13179: pixelout<=1'b1;
13180: pixelout<=1'b1;
13181: pixelout<=1'b1;
13182: pixelout<=1'b1;
13183: pixelout<=1'b1;
13184: pixelout<=1'b1;
13185: pixelout<=1'b1;
13186: pixelout<=1'b1;
13187: pixelout<=1'b1;
13188: pixelout<=1'b1;
13189: pixelout<=1'b1;
13190: pixelout<=1'b1;
13191: pixelout<=1'b1;
13192: pixelout<=1'b1;
13193: pixelout<=1'b1;
13194: pixelout<=1'b1;
13195: pixelout<=1'b1;
13196: pixelout<=1'b1;
13197: pixelout<=1'b1;
13198: pixelout<=1'b1;
13199: pixelout<=1'b1;
13200: pixelout<=1'b1;
13201: pixelout<=1'b1;
13202: pixelout<=1'b1;
13203: pixelout<=1'b1;
13204: pixelout<=1'b1;
13205: pixelout<=1'b1;
13206: pixelout<=1'b1;
13207: pixelout<=1'b1;
13208: pixelout<=1'b1;
13209: pixelout<=1'b1;
13210: pixelout<=1'b1;
13211: pixelout<=1'b1;
13212: pixelout<=1'b1;
13213: pixelout<=1'b1;
13214: pixelout<=1'b1;
13215: pixelout<=1'b1;
13216: pixelout<=1'b1;
13217: pixelout<=1'b1;
13218: pixelout<=1'b1;
13219: pixelout<=1'b1;
13220: pixelout<=1'b1;
13221: pixelout<=1'b1;
13222: pixelout<=1'b1;
13223: pixelout<=1'b1;
13224: pixelout<=1'b1;
13225: pixelout<=1'b1;
13226: pixelout<=1'b1;
13227: pixelout<=1'b1;
13228: pixelout<=1'b1;
13229: pixelout<=1'b1;
13230: pixelout<=1'b1;
13231: pixelout<=1'b1;
13232: pixelout<=1'b0;
13233: pixelout<=1'b1;
13234: pixelout<=1'b1;
13235: pixelout<=1'b1;
13236: pixelout<=1'b1;
13237: pixelout<=1'b1;
13238: pixelout<=1'b1;
13239: pixelout<=1'b1;
13240: pixelout<=1'b0;
13241: pixelout<=1'b1;
13242: pixelout<=1'b0;
13243: pixelout<=1'b1;
13244: pixelout<=1'b1;
13245: pixelout<=1'b1;
13246: pixelout<=1'b0;
13247: pixelout<=1'b1;
13248: pixelout<=1'b0;
13249: pixelout<=1'b1;
13250: pixelout<=1'b1;
13251: pixelout<=1'b1;
13252: pixelout<=1'b0;
13253: pixelout<=1'b1;
13254: pixelout<=1'b0;
13255: pixelout<=1'b1;
13256: pixelout<=1'b0;
13257: pixelout<=1'b1;
13258: pixelout<=1'b1;
13259: pixelout<=1'b1;
13260: pixelout<=1'b1;
13261: pixelout<=1'b1;
13262: pixelout<=1'b1;
13263: pixelout<=1'b1;
13264: pixelout<=1'b1;
13265: pixelout<=1'b1;
13266: pixelout<=1'b1;
13267: pixelout<=1'b1;
13268: pixelout<=1'b1;
13269: pixelout<=1'b0;
13270: pixelout<=1'b1;
13271: pixelout<=1'b1;
13272: pixelout<=1'b1;
13273: pixelout<=1'b0;
13274: pixelout<=1'b1;
13275: pixelout<=1'b1;
13276: pixelout<=1'b1;
13277: pixelout<=1'b0;
13278: pixelout<=1'b1;
13279: pixelout<=1'b0;
13280: pixelout<=1'b1;
13281: pixelout<=1'b1;
13282: pixelout<=1'b1;
13283: pixelout<=1'b1;
13284: pixelout<=1'b1;
13285: pixelout<=1'b1;
13286: pixelout<=1'b1;
13287: pixelout<=1'b1;
13288: pixelout<=1'b1;
13289: pixelout<=1'b0;
13290: pixelout<=1'b1;
13291: pixelout<=1'b0;
13292: pixelout<=1'b1;
13293: pixelout<=1'b0;
13294: pixelout<=1'b1;
13295: pixelout<=1'b1;
13296: pixelout<=1'b0;
13297: pixelout<=1'b1;
13298: pixelout<=1'b1;
13299: pixelout<=1'b1;
13300: pixelout<=1'b1;
13301: pixelout<=1'b1;
13302: pixelout<=1'b1;
13303: pixelout<=1'b1;
13304: pixelout<=1'b0;
13305: pixelout<=1'b1;
13306: pixelout<=1'b1;
13307: pixelout<=1'b1;
13308: pixelout<=1'b0;
13309: pixelout<=1'b1;
13310: pixelout<=1'b1;
13311: pixelout<=1'b1;
13312: pixelout<=1'b1;
13313: pixelout<=1'b1;
13314: pixelout<=1'b1;
13315: pixelout<=1'b1;
13316: pixelout<=1'b1;
13317: pixelout<=1'b0;
13318: pixelout<=1'b1;
13319: pixelout<=1'b1;
13320: pixelout<=1'b1;
13321: pixelout<=1'b0;
13322: pixelout<=1'b1;
13323: pixelout<=1'b0;
13324: pixelout<=1'b1;
13325: pixelout<=1'b1;
13326: pixelout<=1'b0;
13327: pixelout<=1'b1;
13328: pixelout<=1'b1;
13329: pixelout<=1'b0;
13330: pixelout<=1'b0;
13331: pixelout<=1'b1;
13332: pixelout<=1'b1;
13333: pixelout<=1'b1;
13334: pixelout<=1'b1;
13335: pixelout<=1'b1;
13336: pixelout<=1'b1;
13337: pixelout<=1'b1;
13338: pixelout<=1'b1;
13339: pixelout<=1'b0;
13340: pixelout<=1'b1;
13341: pixelout<=1'b1;
13342: pixelout<=1'b1;
13343: pixelout<=1'b0;
13344: pixelout<=1'b0;
13345: pixelout<=1'b0;
13346: pixelout<=1'b0;
13347: pixelout<=1'b0;
13348: pixelout<=1'b1;
13349: pixelout<=1'b1;
13350: pixelout<=1'b1;
13351: pixelout<=1'b0;
13352: pixelout<=1'b1;
13353: pixelout<=1'b1;
13354: pixelout<=1'b1;
13355: pixelout<=1'b0;
13356: pixelout<=1'b1;
13357: pixelout<=1'b0;
13358: pixelout<=1'b1;
13359: pixelout<=1'b1;
13360: pixelout<=1'b1;
13361: pixelout<=1'b1;
13362: pixelout<=1'b1;
13363: pixelout<=1'b1;
13364: pixelout<=1'b1;
13365: pixelout<=1'b1;
13366: pixelout<=1'b1;
13367: pixelout<=1'b1;
13368: pixelout<=1'b0;
13369: pixelout<=1'b1;
13370: pixelout<=1'b0;
13371: pixelout<=1'b1;
13372: pixelout<=1'b1;
13373: pixelout<=1'b0;
13374: pixelout<=1'b1;
13375: pixelout<=1'b1;
13376: pixelout<=1'b0;
13377: pixelout<=1'b1;
13378: pixelout<=1'b1;
13379: pixelout<=1'b0;
13380: pixelout<=1'b1;
13381: pixelout<=1'b1;
13382: pixelout<=1'b1;
13383: pixelout<=1'b1;
13384: pixelout<=1'b1;
13385: pixelout<=1'b1;
13386: pixelout<=1'b1;
13387: pixelout<=1'b1;
13388: pixelout<=1'b1;
13389: pixelout<=1'b1;
13390: pixelout<=1'b1;
13391: pixelout<=1'b1;
13392: pixelout<=1'b1;
13393: pixelout<=1'b1;
13394: pixelout<=1'b0;
13395: pixelout<=1'b1;
13396: pixelout<=1'b0;
13397: pixelout<=1'b1;
13398: pixelout<=1'b1;
13399: pixelout<=1'b1;
13400: pixelout<=1'b0;
13401: pixelout<=1'b1;
13402: pixelout<=1'b0;
13403: pixelout<=1'b1;
13404: pixelout<=1'b1;
13405: pixelout<=1'b0;
13406: pixelout<=1'b1;
13407: pixelout<=1'b1;
13408: pixelout<=1'b1;
13409: pixelout<=1'b1;
13410: pixelout<=1'b1;
13411: pixelout<=1'b1;
13412: pixelout<=1'b1;
13413: pixelout<=1'b1;
13414: pixelout<=1'b1;
13415: pixelout<=1'b1;
13416: pixelout<=1'b1;
13417: pixelout<=1'b1;
13418: pixelout<=1'b1;
13419: pixelout<=1'b1;
13420: pixelout<=1'b1;
13421: pixelout<=1'b1;
13422: pixelout<=1'b1;
13423: pixelout<=1'b1;
13424: pixelout<=1'b1;
13425: pixelout<=1'b1;
13426: pixelout<=1'b1;
13427: pixelout<=1'b1;
13428: pixelout<=1'b1;
13429: pixelout<=1'b1;
13430: pixelout<=1'b1;
13431: pixelout<=1'b1;
13432: pixelout<=1'b1;
13433: pixelout<=1'b1;
13434: pixelout<=1'b1;
13435: pixelout<=1'b1;
13436: pixelout<=1'b1;
13437: pixelout<=1'b1;
13438: pixelout<=1'b1;
13439: pixelout<=1'b1;
13440: pixelout<=1'b1;
13441: pixelout<=1'b1;
13442: pixelout<=1'b1;
13443: pixelout<=1'b1;
13444: pixelout<=1'b1;
13445: pixelout<=1'b1;
13446: pixelout<=1'b1;
13447: pixelout<=1'b1;
13448: pixelout<=1'b1;
13449: pixelout<=1'b1;
13450: pixelout<=1'b1;
13451: pixelout<=1'b1;
13452: pixelout<=1'b1;
13453: pixelout<=1'b1;
13454: pixelout<=1'b1;
13455: pixelout<=1'b1;
13456: pixelout<=1'b1;
13457: pixelout<=1'b1;
13458: pixelout<=1'b1;
13459: pixelout<=1'b1;
13460: pixelout<=1'b1;
13461: pixelout<=1'b1;
13462: pixelout<=1'b1;
13463: pixelout<=1'b1;
13464: pixelout<=1'b1;
13465: pixelout<=1'b1;
13466: pixelout<=1'b1;
13467: pixelout<=1'b1;
13468: pixelout<=1'b1;
13469: pixelout<=1'b1;
13470: pixelout<=1'b1;
13471: pixelout<=1'b1;
13472: pixelout<=1'b1;
13473: pixelout<=1'b1;
13474: pixelout<=1'b1;
13475: pixelout<=1'b1;
13476: pixelout<=1'b1;
13477: pixelout<=1'b1;
13478: pixelout<=1'b1;
13479: pixelout<=1'b1;
13480: pixelout<=1'b0;
13481: pixelout<=1'b1;
13482: pixelout<=1'b0;
13483: pixelout<=1'b0;
13484: pixelout<=1'b0;
13485: pixelout<=1'b0;
13486: pixelout<=1'b0;
13487: pixelout<=1'b1;
13488: pixelout<=1'b0;
13489: pixelout<=1'b1;
13490: pixelout<=1'b1;
13491: pixelout<=1'b1;
13492: pixelout<=1'b1;
13493: pixelout<=1'b1;
13494: pixelout<=1'b0;
13495: pixelout<=1'b1;
13496: pixelout<=1'b0;
13497: pixelout<=1'b1;
13498: pixelout<=1'b1;
13499: pixelout<=1'b1;
13500: pixelout<=1'b1;
13501: pixelout<=1'b1;
13502: pixelout<=1'b1;
13503: pixelout<=1'b1;
13504: pixelout<=1'b1;
13505: pixelout<=1'b1;
13506: pixelout<=1'b1;
13507: pixelout<=1'b1;
13508: pixelout<=1'b1;
13509: pixelout<=1'b0;
13510: pixelout<=1'b1;
13511: pixelout<=1'b1;
13512: pixelout<=1'b1;
13513: pixelout<=1'b0;
13514: pixelout<=1'b1;
13515: pixelout<=1'b1;
13516: pixelout<=1'b1;
13517: pixelout<=1'b0;
13518: pixelout<=1'b1;
13519: pixelout<=1'b0;
13520: pixelout<=1'b1;
13521: pixelout<=1'b1;
13522: pixelout<=1'b1;
13523: pixelout<=1'b1;
13524: pixelout<=1'b1;
13525: pixelout<=1'b1;
13526: pixelout<=1'b1;
13527: pixelout<=1'b1;
13528: pixelout<=1'b1;
13529: pixelout<=1'b0;
13530: pixelout<=1'b1;
13531: pixelout<=1'b0;
13532: pixelout<=1'b0;
13533: pixelout<=1'b1;
13534: pixelout<=1'b1;
13535: pixelout<=1'b1;
13536: pixelout<=1'b1;
13537: pixelout<=1'b0;
13538: pixelout<=1'b0;
13539: pixelout<=1'b1;
13540: pixelout<=1'b1;
13541: pixelout<=1'b1;
13542: pixelout<=1'b1;
13543: pixelout<=1'b1;
13544: pixelout<=1'b0;
13545: pixelout<=1'b1;
13546: pixelout<=1'b1;
13547: pixelout<=1'b1;
13548: pixelout<=1'b0;
13549: pixelout<=1'b1;
13550: pixelout<=1'b1;
13551: pixelout<=1'b1;
13552: pixelout<=1'b1;
13553: pixelout<=1'b1;
13554: pixelout<=1'b1;
13555: pixelout<=1'b1;
13556: pixelout<=1'b1;
13557: pixelout<=1'b0;
13558: pixelout<=1'b1;
13559: pixelout<=1'b1;
13560: pixelout<=1'b1;
13561: pixelout<=1'b0;
13562: pixelout<=1'b1;
13563: pixelout<=1'b0;
13564: pixelout<=1'b1;
13565: pixelout<=1'b1;
13566: pixelout<=1'b0;
13567: pixelout<=1'b1;
13568: pixelout<=1'b1;
13569: pixelout<=1'b0;
13570: pixelout<=1'b1;
13571: pixelout<=1'b1;
13572: pixelout<=1'b1;
13573: pixelout<=1'b1;
13574: pixelout<=1'b1;
13575: pixelout<=1'b1;
13576: pixelout<=1'b1;
13577: pixelout<=1'b1;
13578: pixelout<=1'b1;
13579: pixelout<=1'b0;
13580: pixelout<=1'b1;
13581: pixelout<=1'b1;
13582: pixelout<=1'b1;
13583: pixelout<=1'b0;
13584: pixelout<=1'b1;
13585: pixelout<=1'b1;
13586: pixelout<=1'b1;
13587: pixelout<=1'b0;
13588: pixelout<=1'b1;
13589: pixelout<=1'b1;
13590: pixelout<=1'b1;
13591: pixelout<=1'b0;
13592: pixelout<=1'b1;
13593: pixelout<=1'b1;
13594: pixelout<=1'b1;
13595: pixelout<=1'b0;
13596: pixelout<=1'b1;
13597: pixelout<=1'b0;
13598: pixelout<=1'b1;
13599: pixelout<=1'b1;
13600: pixelout<=1'b1;
13601: pixelout<=1'b1;
13602: pixelout<=1'b1;
13603: pixelout<=1'b1;
13604: pixelout<=1'b1;
13605: pixelout<=1'b1;
13606: pixelout<=1'b1;
13607: pixelout<=1'b1;
13608: pixelout<=1'b0;
13609: pixelout<=1'b1;
13610: pixelout<=1'b0;
13611: pixelout<=1'b1;
13612: pixelout<=1'b1;
13613: pixelout<=1'b0;
13614: pixelout<=1'b1;
13615: pixelout<=1'b1;
13616: pixelout<=1'b0;
13617: pixelout<=1'b1;
13618: pixelout<=1'b1;
13619: pixelout<=1'b0;
13620: pixelout<=1'b1;
13621: pixelout<=1'b1;
13622: pixelout<=1'b1;
13623: pixelout<=1'b1;
13624: pixelout<=1'b1;
13625: pixelout<=1'b1;
13626: pixelout<=1'b1;
13627: pixelout<=1'b1;
13628: pixelout<=1'b1;
13629: pixelout<=1'b1;
13630: pixelout<=1'b0;
13631: pixelout<=1'b0;
13632: pixelout<=1'b0;
13633: pixelout<=1'b0;
13634: pixelout<=1'b0;
13635: pixelout<=1'b1;
13636: pixelout<=1'b0;
13637: pixelout<=1'b1;
13638: pixelout<=1'b1;
13639: pixelout<=1'b1;
13640: pixelout<=1'b0;
13641: pixelout<=1'b1;
13642: pixelout<=1'b0;
13643: pixelout<=1'b1;
13644: pixelout<=1'b1;
13645: pixelout<=1'b0;
13646: pixelout<=1'b1;
13647: pixelout<=1'b1;
13648: pixelout<=1'b1;
13649: pixelout<=1'b1;
13650: pixelout<=1'b1;
13651: pixelout<=1'b1;
13652: pixelout<=1'b1;
13653: pixelout<=1'b1;
13654: pixelout<=1'b1;
13655: pixelout<=1'b1;
13656: pixelout<=1'b1;
13657: pixelout<=1'b1;
13658: pixelout<=1'b1;
13659: pixelout<=1'b1;
13660: pixelout<=1'b1;
13661: pixelout<=1'b1;
13662: pixelout<=1'b1;
13663: pixelout<=1'b1;
13664: pixelout<=1'b1;
13665: pixelout<=1'b1;
13666: pixelout<=1'b1;
13667: pixelout<=1'b1;
13668: pixelout<=1'b1;
13669: pixelout<=1'b1;
13670: pixelout<=1'b1;
13671: pixelout<=1'b1;
13672: pixelout<=1'b1;
13673: pixelout<=1'b1;
13674: pixelout<=1'b1;
13675: pixelout<=1'b1;
13676: pixelout<=1'b1;
13677: pixelout<=1'b1;
13678: pixelout<=1'b1;
13679: pixelout<=1'b1;
13680: pixelout<=1'b1;
13681: pixelout<=1'b1;
13682: pixelout<=1'b1;
13683: pixelout<=1'b1;
13684: pixelout<=1'b1;
13685: pixelout<=1'b1;
13686: pixelout<=1'b1;
13687: pixelout<=1'b1;
13688: pixelout<=1'b1;
13689: pixelout<=1'b1;
13690: pixelout<=1'b1;
13691: pixelout<=1'b1;
13692: pixelout<=1'b1;
13693: pixelout<=1'b1;
13694: pixelout<=1'b1;
13695: pixelout<=1'b1;
13696: pixelout<=1'b1;
13697: pixelout<=1'b1;
13698: pixelout<=1'b1;
13699: pixelout<=1'b1;
13700: pixelout<=1'b1;
13701: pixelout<=1'b1;
13702: pixelout<=1'b1;
13703: pixelout<=1'b1;
13704: pixelout<=1'b1;
13705: pixelout<=1'b1;
13706: pixelout<=1'b1;
13707: pixelout<=1'b1;
13708: pixelout<=1'b1;
13709: pixelout<=1'b0;
13710: pixelout<=1'b1;
13711: pixelout<=1'b1;
13712: pixelout<=1'b1;
13713: pixelout<=1'b1;
13714: pixelout<=1'b1;
13715: pixelout<=1'b1;
13716: pixelout<=1'b1;
13717: pixelout<=1'b1;
13718: pixelout<=1'b1;
13719: pixelout<=1'b1;
13720: pixelout<=1'b0;
13721: pixelout<=1'b1;
13722: pixelout<=1'b0;
13723: pixelout<=1'b1;
13724: pixelout<=1'b1;
13725: pixelout<=1'b1;
13726: pixelout<=1'b1;
13727: pixelout<=1'b1;
13728: pixelout<=1'b0;
13729: pixelout<=1'b1;
13730: pixelout<=1'b1;
13731: pixelout<=1'b1;
13732: pixelout<=1'b0;
13733: pixelout<=1'b1;
13734: pixelout<=1'b0;
13735: pixelout<=1'b1;
13736: pixelout<=1'b0;
13737: pixelout<=1'b1;
13738: pixelout<=1'b1;
13739: pixelout<=1'b0;
13740: pixelout<=1'b0;
13741: pixelout<=1'b1;
13742: pixelout<=1'b1;
13743: pixelout<=1'b1;
13744: pixelout<=1'b1;
13745: pixelout<=1'b1;
13746: pixelout<=1'b1;
13747: pixelout<=1'b1;
13748: pixelout<=1'b1;
13749: pixelout<=1'b0;
13750: pixelout<=1'b1;
13751: pixelout<=1'b1;
13752: pixelout<=1'b1;
13753: pixelout<=1'b0;
13754: pixelout<=1'b1;
13755: pixelout<=1'b1;
13756: pixelout<=1'b1;
13757: pixelout<=1'b0;
13758: pixelout<=1'b1;
13759: pixelout<=1'b0;
13760: pixelout<=1'b1;
13761: pixelout<=1'b1;
13762: pixelout<=1'b0;
13763: pixelout<=1'b0;
13764: pixelout<=1'b1;
13765: pixelout<=1'b1;
13766: pixelout<=1'b1;
13767: pixelout<=1'b1;
13768: pixelout<=1'b1;
13769: pixelout<=1'b0;
13770: pixelout<=1'b1;
13771: pixelout<=1'b0;
13772: pixelout<=1'b1;
13773: pixelout<=1'b0;
13774: pixelout<=1'b1;
13775: pixelout<=1'b1;
13776: pixelout<=1'b1;
13777: pixelout<=1'b1;
13778: pixelout<=1'b1;
13779: pixelout<=1'b0;
13780: pixelout<=1'b1;
13781: pixelout<=1'b1;
13782: pixelout<=1'b1;
13783: pixelout<=1'b1;
13784: pixelout<=1'b0;
13785: pixelout<=1'b1;
13786: pixelout<=1'b1;
13787: pixelout<=1'b1;
13788: pixelout<=1'b0;
13789: pixelout<=1'b1;
13790: pixelout<=1'b1;
13791: pixelout<=1'b1;
13792: pixelout<=1'b1;
13793: pixelout<=1'b1;
13794: pixelout<=1'b1;
13795: pixelout<=1'b1;
13796: pixelout<=1'b1;
13797: pixelout<=1'b0;
13798: pixelout<=1'b1;
13799: pixelout<=1'b1;
13800: pixelout<=1'b1;
13801: pixelout<=1'b0;
13802: pixelout<=1'b1;
13803: pixelout<=1'b0;
13804: pixelout<=1'b1;
13805: pixelout<=1'b1;
13806: pixelout<=1'b0;
13807: pixelout<=1'b1;
13808: pixelout<=1'b1;
13809: pixelout<=1'b0;
13810: pixelout<=1'b1;
13811: pixelout<=1'b1;
13812: pixelout<=1'b1;
13813: pixelout<=1'b1;
13814: pixelout<=1'b1;
13815: pixelout<=1'b1;
13816: pixelout<=1'b1;
13817: pixelout<=1'b1;
13818: pixelout<=1'b1;
13819: pixelout<=1'b0;
13820: pixelout<=1'b1;
13821: pixelout<=1'b1;
13822: pixelout<=1'b1;
13823: pixelout<=1'b0;
13824: pixelout<=1'b1;
13825: pixelout<=1'b1;
13826: pixelout<=1'b1;
13827: pixelout<=1'b0;
13828: pixelout<=1'b1;
13829: pixelout<=1'b1;
13830: pixelout<=1'b1;
13831: pixelout<=1'b0;
13832: pixelout<=1'b1;
13833: pixelout<=1'b1;
13834: pixelout<=1'b1;
13835: pixelout<=1'b0;
13836: pixelout<=1'b1;
13837: pixelout<=1'b0;
13838: pixelout<=1'b1;
13839: pixelout<=1'b1;
13840: pixelout<=1'b1;
13841: pixelout<=1'b1;
13842: pixelout<=1'b1;
13843: pixelout<=1'b1;
13844: pixelout<=1'b1;
13845: pixelout<=1'b1;
13846: pixelout<=1'b1;
13847: pixelout<=1'b1;
13848: pixelout<=1'b0;
13849: pixelout<=1'b1;
13850: pixelout<=1'b0;
13851: pixelout<=1'b1;
13852: pixelout<=1'b1;
13853: pixelout<=1'b0;
13854: pixelout<=1'b1;
13855: pixelout<=1'b1;
13856: pixelout<=1'b0;
13857: pixelout<=1'b1;
13858: pixelout<=1'b1;
13859: pixelout<=1'b0;
13860: pixelout<=1'b1;
13861: pixelout<=1'b1;
13862: pixelout<=1'b1;
13863: pixelout<=1'b0;
13864: pixelout<=1'b1;
13865: pixelout<=1'b1;
13866: pixelout<=1'b1;
13867: pixelout<=1'b1;
13868: pixelout<=1'b1;
13869: pixelout<=1'b1;
13870: pixelout<=1'b1;
13871: pixelout<=1'b1;
13872: pixelout<=1'b1;
13873: pixelout<=1'b1;
13874: pixelout<=1'b1;
13875: pixelout<=1'b1;
13876: pixelout<=1'b0;
13877: pixelout<=1'b1;
13878: pixelout<=1'b1;
13879: pixelout<=1'b1;
13880: pixelout<=1'b0;
13881: pixelout<=1'b1;
13882: pixelout<=1'b0;
13883: pixelout<=1'b1;
13884: pixelout<=1'b1;
13885: pixelout<=1'b0;
13886: pixelout<=1'b1;
13887: pixelout<=1'b0;
13888: pixelout<=1'b0;
13889: pixelout<=1'b1;
13890: pixelout<=1'b1;
13891: pixelout<=1'b1;
13892: pixelout<=1'b1;
13893: pixelout<=1'b1;
13894: pixelout<=1'b1;
13895: pixelout<=1'b1;
13896: pixelout<=1'b1;
13897: pixelout<=1'b1;
13898: pixelout<=1'b1;
13899: pixelout<=1'b1;
13900: pixelout<=1'b1;
13901: pixelout<=1'b1;
13902: pixelout<=1'b1;
13903: pixelout<=1'b1;
13904: pixelout<=1'b1;
13905: pixelout<=1'b1;
13906: pixelout<=1'b1;
13907: pixelout<=1'b1;
13908: pixelout<=1'b1;
13909: pixelout<=1'b1;
13910: pixelout<=1'b1;
13911: pixelout<=1'b1;
13912: pixelout<=1'b1;
13913: pixelout<=1'b1;
13914: pixelout<=1'b1;
13915: pixelout<=1'b1;
13916: pixelout<=1'b1;
13917: pixelout<=1'b1;
13918: pixelout<=1'b1;
13919: pixelout<=1'b1;
13920: pixelout<=1'b1;
13921: pixelout<=1'b1;
13922: pixelout<=1'b1;
13923: pixelout<=1'b1;
13924: pixelout<=1'b1;
13925: pixelout<=1'b1;
13926: pixelout<=1'b1;
13927: pixelout<=1'b1;
13928: pixelout<=1'b1;
13929: pixelout<=1'b1;
13930: pixelout<=1'b1;
13931: pixelout<=1'b1;
13932: pixelout<=1'b1;
13933: pixelout<=1'b1;
13934: pixelout<=1'b1;
13935: pixelout<=1'b1;
13936: pixelout<=1'b1;
13937: pixelout<=1'b1;
13938: pixelout<=1'b1;
13939: pixelout<=1'b1;
13940: pixelout<=1'b1;
13941: pixelout<=1'b1;
13942: pixelout<=1'b1;
13943: pixelout<=1'b1;
13944: pixelout<=1'b1;
13945: pixelout<=1'b1;
13946: pixelout<=1'b1;
13947: pixelout<=1'b1;
13948: pixelout<=1'b1;
13949: pixelout<=1'b1;
13950: pixelout<=1'b0;
13951: pixelout<=1'b0;
13952: pixelout<=1'b0;
13953: pixelout<=1'b1;
13954: pixelout<=1'b1;
13955: pixelout<=1'b1;
13956: pixelout<=1'b0;
13957: pixelout<=1'b0;
13958: pixelout<=1'b0;
13959: pixelout<=1'b0;
13960: pixelout<=1'b1;
13961: pixelout<=1'b1;
13962: pixelout<=1'b1;
13963: pixelout<=1'b0;
13964: pixelout<=1'b0;
13965: pixelout<=1'b0;
13966: pixelout<=1'b0;
13967: pixelout<=1'b1;
13968: pixelout<=1'b1;
13969: pixelout<=1'b0;
13970: pixelout<=1'b0;
13971: pixelout<=1'b0;
13972: pixelout<=1'b1;
13973: pixelout<=1'b1;
13974: pixelout<=1'b0;
13975: pixelout<=1'b1;
13976: pixelout<=1'b1;
13977: pixelout<=1'b0;
13978: pixelout<=1'b0;
13979: pixelout<=1'b1;
13980: pixelout<=1'b1;
13981: pixelout<=1'b1;
13982: pixelout<=1'b1;
13983: pixelout<=1'b1;
13984: pixelout<=1'b1;
13985: pixelout<=1'b1;
13986: pixelout<=1'b1;
13987: pixelout<=1'b1;
13988: pixelout<=1'b1;
13989: pixelout<=1'b0;
13990: pixelout<=1'b0;
13991: pixelout<=1'b0;
13992: pixelout<=1'b1;
13993: pixelout<=1'b0;
13994: pixelout<=1'b1;
13995: pixelout<=1'b1;
13996: pixelout<=1'b1;
13997: pixelout<=1'b0;
13998: pixelout<=1'b1;
13999: pixelout<=1'b1;
14000: pixelout<=1'b0;
14001: pixelout<=1'b0;
14002: pixelout<=1'b1;
14003: pixelout<=1'b1;
14004: pixelout<=1'b1;
14005: pixelout<=1'b1;
14006: pixelout<=1'b1;
14007: pixelout<=1'b1;
14008: pixelout<=1'b1;
14009: pixelout<=1'b0;
14010: pixelout<=1'b1;
14011: pixelout<=1'b0;
14012: pixelout<=1'b1;
14013: pixelout<=1'b1;
14014: pixelout<=1'b0;
14015: pixelout<=1'b1;
14016: pixelout<=1'b0;
14017: pixelout<=1'b0;
14018: pixelout<=1'b0;
14019: pixelout<=1'b0;
14020: pixelout<=1'b1;
14021: pixelout<=1'b1;
14022: pixelout<=1'b1;
14023: pixelout<=1'b1;
14024: pixelout<=1'b0;
14025: pixelout<=1'b0;
14026: pixelout<=1'b0;
14027: pixelout<=1'b1;
14028: pixelout<=1'b1;
14029: pixelout<=1'b0;
14030: pixelout<=1'b0;
14031: pixelout<=1'b0;
14032: pixelout<=1'b1;
14033: pixelout<=1'b1;
14034: pixelout<=1'b1;
14035: pixelout<=1'b1;
14036: pixelout<=1'b1;
14037: pixelout<=1'b1;
14038: pixelout<=1'b0;
14039: pixelout<=1'b0;
14040: pixelout<=1'b0;
14041: pixelout<=1'b1;
14042: pixelout<=1'b1;
14043: pixelout<=1'b1;
14044: pixelout<=1'b0;
14045: pixelout<=1'b0;
14046: pixelout<=1'b1;
14047: pixelout<=1'b0;
14048: pixelout<=1'b1;
14049: pixelout<=1'b0;
14050: pixelout<=1'b1;
14051: pixelout<=1'b1;
14052: pixelout<=1'b1;
14053: pixelout<=1'b1;
14054: pixelout<=1'b1;
14055: pixelout<=1'b1;
14056: pixelout<=1'b1;
14057: pixelout<=1'b1;
14058: pixelout<=1'b1;
14059: pixelout<=1'b0;
14060: pixelout<=1'b1;
14061: pixelout<=1'b1;
14062: pixelout<=1'b1;
14063: pixelout<=1'b0;
14064: pixelout<=1'b1;
14065: pixelout<=1'b1;
14066: pixelout<=1'b1;
14067: pixelout<=1'b0;
14068: pixelout<=1'b1;
14069: pixelout<=1'b1;
14070: pixelout<=1'b1;
14071: pixelout<=1'b0;
14072: pixelout<=1'b0;
14073: pixelout<=1'b0;
14074: pixelout<=1'b0;
14075: pixelout<=1'b1;
14076: pixelout<=1'b1;
14077: pixelout<=1'b1;
14078: pixelout<=1'b0;
14079: pixelout<=1'b0;
14080: pixelout<=1'b0;
14081: pixelout<=1'b1;
14082: pixelout<=1'b1;
14083: pixelout<=1'b1;
14084: pixelout<=1'b1;
14085: pixelout<=1'b1;
14086: pixelout<=1'b1;
14087: pixelout<=1'b1;
14088: pixelout<=1'b0;
14089: pixelout<=1'b1;
14090: pixelout<=1'b1;
14091: pixelout<=1'b0;
14092: pixelout<=1'b0;
14093: pixelout<=1'b1;
14094: pixelout<=1'b0;
14095: pixelout<=1'b1;
14096: pixelout<=1'b0;
14097: pixelout<=1'b1;
14098: pixelout<=1'b1;
14099: pixelout<=1'b0;
14100: pixelout<=1'b1;
14101: pixelout<=1'b1;
14102: pixelout<=1'b1;
14103: pixelout<=1'b1;
14104: pixelout<=1'b0;
14105: pixelout<=1'b0;
14106: pixelout<=1'b0;
14107: pixelout<=1'b1;
14108: pixelout<=1'b1;
14109: pixelout<=1'b1;
14110: pixelout<=1'b1;
14111: pixelout<=1'b0;
14112: pixelout<=1'b0;
14113: pixelout<=1'b0;
14114: pixelout<=1'b0;
14115: pixelout<=1'b1;
14116: pixelout<=1'b1;
14117: pixelout<=1'b0;
14118: pixelout<=1'b0;
14119: pixelout<=1'b0;
14120: pixelout<=1'b1;
14121: pixelout<=1'b1;
14122: pixelout<=1'b0;
14123: pixelout<=1'b1;
14124: pixelout<=1'b1;
14125: pixelout<=1'b0;
14126: pixelout<=1'b1;
14127: pixelout<=1'b0;
14128: pixelout<=1'b0;
14129: pixelout<=1'b1;
14130: pixelout<=1'b1;
14131: pixelout<=1'b1;
14132: pixelout<=1'b1;
14133: pixelout<=1'b1;
14134: pixelout<=1'b1;
14135: pixelout<=1'b1;
14136: pixelout<=1'b1;
14137: pixelout<=1'b1;
14138: pixelout<=1'b1;
14139: pixelout<=1'b1;
14140: pixelout<=1'b1;
14141: pixelout<=1'b1;
14142: pixelout<=1'b1;
14143: pixelout<=1'b1;
14144: pixelout<=1'b1;
14145: pixelout<=1'b1;
14146: pixelout<=1'b1;
14147: pixelout<=1'b1;
14148: pixelout<=1'b1;
14149: pixelout<=1'b1;
14150: pixelout<=1'b1;
14151: pixelout<=1'b1;
14152: pixelout<=1'b1;
14153: pixelout<=1'b1;
14154: pixelout<=1'b1;
14155: pixelout<=1'b1;
14156: pixelout<=1'b1;
14157: pixelout<=1'b1;
14158: pixelout<=1'b1;
14159: pixelout<=1'b1;
14160: pixelout<=1'b1;
14161: pixelout<=1'b1;
14162: pixelout<=1'b1;
14163: pixelout<=1'b1;
14164: pixelout<=1'b1;
14165: pixelout<=1'b1;
14166: pixelout<=1'b1;
14167: pixelout<=1'b1;
14168: pixelout<=1'b1;
14169: pixelout<=1'b1;
14170: pixelout<=1'b1;
14171: pixelout<=1'b1;
14172: pixelout<=1'b1;
14173: pixelout<=1'b1;
14174: pixelout<=1'b1;
14175: pixelout<=1'b1;
14176: pixelout<=1'b1;
14177: pixelout<=1'b1;
14178: pixelout<=1'b1;
14179: pixelout<=1'b1;
14180: pixelout<=1'b1;
14181: pixelout<=1'b1;
14182: pixelout<=1'b1;
14183: pixelout<=1'b1;
14184: pixelout<=1'b1;
14185: pixelout<=1'b1;
14186: pixelout<=1'b1;
14187: pixelout<=1'b1;
14188: pixelout<=1'b1;
14189: pixelout<=1'b1;
14190: pixelout<=1'b1;
14191: pixelout<=1'b1;
14192: pixelout<=1'b1;
14193: pixelout<=1'b1;
14194: pixelout<=1'b1;
14195: pixelout<=1'b1;
14196: pixelout<=1'b1;
14197: pixelout<=1'b1;
14198: pixelout<=1'b1;
14199: pixelout<=1'b1;
14200: pixelout<=1'b1;
14201: pixelout<=1'b1;
14202: pixelout<=1'b1;
14203: pixelout<=1'b1;
14204: pixelout<=1'b1;
14205: pixelout<=1'b1;
14206: pixelout<=1'b1;
14207: pixelout<=1'b1;
14208: pixelout<=1'b1;
14209: pixelout<=1'b1;
14210: pixelout<=1'b1;
14211: pixelout<=1'b1;
14212: pixelout<=1'b1;
14213: pixelout<=1'b1;
14214: pixelout<=1'b1;
14215: pixelout<=1'b1;
14216: pixelout<=1'b1;
14217: pixelout<=1'b1;
14218: pixelout<=1'b1;
14219: pixelout<=1'b1;
14220: pixelout<=1'b1;
14221: pixelout<=1'b1;
14222: pixelout<=1'b1;
14223: pixelout<=1'b1;
14224: pixelout<=1'b1;
14225: pixelout<=1'b1;
14226: pixelout<=1'b1;
14227: pixelout<=1'b1;
14228: pixelout<=1'b1;
14229: pixelout<=1'b1;
14230: pixelout<=1'b1;
14231: pixelout<=1'b1;
14232: pixelout<=1'b1;
14233: pixelout<=1'b1;
14234: pixelout<=1'b1;
14235: pixelout<=1'b1;
14236: pixelout<=1'b1;
14237: pixelout<=1'b1;
14238: pixelout<=1'b1;
14239: pixelout<=1'b1;
14240: pixelout<=1'b1;
14241: pixelout<=1'b1;
14242: pixelout<=1'b1;
14243: pixelout<=1'b1;
14244: pixelout<=1'b1;
14245: pixelout<=1'b1;
14246: pixelout<=1'b1;
14247: pixelout<=1'b1;
14248: pixelout<=1'b1;
14249: pixelout<=1'b1;
14250: pixelout<=1'b1;
14251: pixelout<=1'b1;
14252: pixelout<=1'b1;
14253: pixelout<=1'b1;
14254: pixelout<=1'b1;
14255: pixelout<=1'b1;
14256: pixelout<=1'b1;
14257: pixelout<=1'b1;
14258: pixelout<=1'b1;
14259: pixelout<=1'b1;
14260: pixelout<=1'b1;
14261: pixelout<=1'b1;
14262: pixelout<=1'b1;
14263: pixelout<=1'b1;
14264: pixelout<=1'b1;
14265: pixelout<=1'b1;
14266: pixelout<=1'b1;
14267: pixelout<=1'b1;
14268: pixelout<=1'b1;
14269: pixelout<=1'b1;
14270: pixelout<=1'b1;
14271: pixelout<=1'b1;
14272: pixelout<=1'b1;
14273: pixelout<=1'b1;
14274: pixelout<=1'b1;
14275: pixelout<=1'b1;
14276: pixelout<=1'b1;
14277: pixelout<=1'b1;
14278: pixelout<=1'b1;
14279: pixelout<=1'b1;
14280: pixelout<=1'b1;
14281: pixelout<=1'b1;
14282: pixelout<=1'b1;
14283: pixelout<=1'b1;
14284: pixelout<=1'b1;
14285: pixelout<=1'b1;
14286: pixelout<=1'b1;
14287: pixelout<=1'b1;
14288: pixelout<=1'b1;
14289: pixelout<=1'b1;
14290: pixelout<=1'b1;
14291: pixelout<=1'b1;
14292: pixelout<=1'b1;
14293: pixelout<=1'b1;
14294: pixelout<=1'b1;
14295: pixelout<=1'b1;
14296: pixelout<=1'b1;
14297: pixelout<=1'b1;
14298: pixelout<=1'b1;
14299: pixelout<=1'b1;
14300: pixelout<=1'b1;
14301: pixelout<=1'b1;
14302: pixelout<=1'b1;
14303: pixelout<=1'b1;
14304: pixelout<=1'b1;
14305: pixelout<=1'b1;
14306: pixelout<=1'b1;
14307: pixelout<=1'b1;
14308: pixelout<=1'b1;
14309: pixelout<=1'b1;
14310: pixelout<=1'b1;
14311: pixelout<=1'b1;
14312: pixelout<=1'b1;
14313: pixelout<=1'b1;
14314: pixelout<=1'b1;
14315: pixelout<=1'b1;
14316: pixelout<=1'b1;
14317: pixelout<=1'b1;
14318: pixelout<=1'b1;
14319: pixelout<=1'b1;
14320: pixelout<=1'b1;
14321: pixelout<=1'b1;
14322: pixelout<=1'b1;
14323: pixelout<=1'b1;
14324: pixelout<=1'b1;
14325: pixelout<=1'b1;
14326: pixelout<=1'b1;
14327: pixelout<=1'b1;
14328: pixelout<=1'b1;
14329: pixelout<=1'b1;
14330: pixelout<=1'b1;
14331: pixelout<=1'b1;
14332: pixelout<=1'b1;
14333: pixelout<=1'b1;
14334: pixelout<=1'b1;
14335: pixelout<=1'b1;
14336: pixelout<=1'b1;
14337: pixelout<=1'b1;
14338: pixelout<=1'b1;
14339: pixelout<=1'b1;
14340: pixelout<=1'b1;
14341: pixelout<=1'b1;
14342: pixelout<=1'b1;
14343: pixelout<=1'b1;
14344: pixelout<=1'b1;
14345: pixelout<=1'b1;
14346: pixelout<=1'b1;
14347: pixelout<=1'b1;
14348: pixelout<=1'b1;
14349: pixelout<=1'b1;
14350: pixelout<=1'b1;
14351: pixelout<=1'b1;
14352: pixelout<=1'b1;
14353: pixelout<=1'b1;
14354: pixelout<=1'b1;
14355: pixelout<=1'b1;
14356: pixelout<=1'b1;
14357: pixelout<=1'b1;
14358: pixelout<=1'b1;
14359: pixelout<=1'b1;
14360: pixelout<=1'b1;
14361: pixelout<=1'b1;
14362: pixelout<=1'b1;
14363: pixelout<=1'b1;
14364: pixelout<=1'b1;
14365: pixelout<=1'b1;
14366: pixelout<=1'b1;
14367: pixelout<=1'b1;
14368: pixelout<=1'b0;
14369: pixelout<=1'b1;
14370: pixelout<=1'b1;
14371: pixelout<=1'b1;
14372: pixelout<=1'b1;
14373: pixelout<=1'b1;
14374: pixelout<=1'b1;
14375: pixelout<=1'b1;
14376: pixelout<=1'b1;
14377: pixelout<=1'b1;
14378: pixelout<=1'b1;
14379: pixelout<=1'b1;
14380: pixelout<=1'b1;
14381: pixelout<=1'b1;
14382: pixelout<=1'b1;
14383: pixelout<=1'b1;
14384: pixelout<=1'b1;
14385: pixelout<=1'b1;
14386: pixelout<=1'b1;
14387: pixelout<=1'b1;
14388: pixelout<=1'b1;
14389: pixelout<=1'b1;
14390: pixelout<=1'b1;
14391: pixelout<=1'b1;
14392: pixelout<=1'b1;
14393: pixelout<=1'b1;
14394: pixelout<=1'b1;
14395: pixelout<=1'b1;
14396: pixelout<=1'b1;
14397: pixelout<=1'b1;
14398: pixelout<=1'b1;
14399: pixelout<=1'b1;
14400: pixelout<=1'b1;
14401: pixelout<=1'b1;
14402: pixelout<=1'b1;
14403: pixelout<=1'b1;
14404: pixelout<=1'b1;
14405: pixelout<=1'b1;
14406: pixelout<=1'b1;
14407: pixelout<=1'b1;
14408: pixelout<=1'b1;
14409: pixelout<=1'b1;
14410: pixelout<=1'b1;
14411: pixelout<=1'b1;
14412: pixelout<=1'b1;
14413: pixelout<=1'b1;
14414: pixelout<=1'b1;
14415: pixelout<=1'b1;
14416: pixelout<=1'b1;
14417: pixelout<=1'b1;
14418: pixelout<=1'b1;
14419: pixelout<=1'b1;
14420: pixelout<=1'b1;
14421: pixelout<=1'b1;
14422: pixelout<=1'b1;
14423: pixelout<=1'b1;
14424: pixelout<=1'b1;
14425: pixelout<=1'b1;
14426: pixelout<=1'b1;
14427: pixelout<=1'b1;
14428: pixelout<=1'b1;
14429: pixelout<=1'b1;
14430: pixelout<=1'b1;
14431: pixelout<=1'b1;
14432: pixelout<=1'b1;
14433: pixelout<=1'b1;
14434: pixelout<=1'b1;
14435: pixelout<=1'b1;
14436: pixelout<=1'b1;
14437: pixelout<=1'b1;
14438: pixelout<=1'b1;
14439: pixelout<=1'b1;
14440: pixelout<=1'b1;
14441: pixelout<=1'b1;
14442: pixelout<=1'b1;
14443: pixelout<=1'b1;
14444: pixelout<=1'b1;
14445: pixelout<=1'b1;
14446: pixelout<=1'b1;
14447: pixelout<=1'b1;
14448: pixelout<=1'b1;
14449: pixelout<=1'b1;
14450: pixelout<=1'b1;
14451: pixelout<=1'b1;
14452: pixelout<=1'b1;
14453: pixelout<=1'b1;
14454: pixelout<=1'b1;
14455: pixelout<=1'b1;
14456: pixelout<=1'b1;
14457: pixelout<=1'b1;
14458: pixelout<=1'b1;
14459: pixelout<=1'b1;
14460: pixelout<=1'b1;
14461: pixelout<=1'b1;
14462: pixelout<=1'b1;
14463: pixelout<=1'b1;
14464: pixelout<=1'b1;
14465: pixelout<=1'b1;
14466: pixelout<=1'b1;
14467: pixelout<=1'b1;
14468: pixelout<=1'b1;
14469: pixelout<=1'b1;
14470: pixelout<=1'b1;
14471: pixelout<=1'b1;
14472: pixelout<=1'b1;
14473: pixelout<=1'b1;
14474: pixelout<=1'b1;
14475: pixelout<=1'b1;
14476: pixelout<=1'b1;
14477: pixelout<=1'b1;
14478: pixelout<=1'b1;
14479: pixelout<=1'b1;
14480: pixelout<=1'b1;
14481: pixelout<=1'b1;
14482: pixelout<=1'b1;
14483: pixelout<=1'b1;
14484: pixelout<=1'b1;
14485: pixelout<=1'b1;
14486: pixelout<=1'b1;
14487: pixelout<=1'b1;
14488: pixelout<=1'b1;
14489: pixelout<=1'b1;
14490: pixelout<=1'b1;
14491: pixelout<=1'b1;
14492: pixelout<=1'b1;
14493: pixelout<=1'b1;
14494: pixelout<=1'b1;
14495: pixelout<=1'b1;
14496: pixelout<=1'b1;
14497: pixelout<=1'b1;
14498: pixelout<=1'b1;
14499: pixelout<=1'b1;
14500: pixelout<=1'b1;
14501: pixelout<=1'b1;
14502: pixelout<=1'b1;
14503: pixelout<=1'b1;
14504: pixelout<=1'b1;
14505: pixelout<=1'b1;
14506: pixelout<=1'b1;
14507: pixelout<=1'b1;
14508: pixelout<=1'b1;
14509: pixelout<=1'b1;
14510: pixelout<=1'b1;
14511: pixelout<=1'b1;
14512: pixelout<=1'b1;
14513: pixelout<=1'b1;
14514: pixelout<=1'b1;
14515: pixelout<=1'b1;
14516: pixelout<=1'b1;
14517: pixelout<=1'b1;
14518: pixelout<=1'b1;
14519: pixelout<=1'b1;
14520: pixelout<=1'b1;
14521: pixelout<=1'b1;
14522: pixelout<=1'b1;
14523: pixelout<=1'b1;
14524: pixelout<=1'b1;
14525: pixelout<=1'b1;
14526: pixelout<=1'b1;
14527: pixelout<=1'b1;
14528: pixelout<=1'b1;
14529: pixelout<=1'b1;
14530: pixelout<=1'b1;
14531: pixelout<=1'b1;
14532: pixelout<=1'b1;
14533: pixelout<=1'b1;
14534: pixelout<=1'b1;
14535: pixelout<=1'b1;
14536: pixelout<=1'b1;
14537: pixelout<=1'b1;
14538: pixelout<=1'b1;
14539: pixelout<=1'b1;
14540: pixelout<=1'b1;
14541: pixelout<=1'b1;
14542: pixelout<=1'b1;
14543: pixelout<=1'b1;
14544: pixelout<=1'b1;
14545: pixelout<=1'b1;
14546: pixelout<=1'b1;
14547: pixelout<=1'b1;
14548: pixelout<=1'b1;
14549: pixelout<=1'b1;
14550: pixelout<=1'b1;
14551: pixelout<=1'b1;
14552: pixelout<=1'b1;
14553: pixelout<=1'b1;
14554: pixelout<=1'b1;
14555: pixelout<=1'b1;
14556: pixelout<=1'b1;
14557: pixelout<=1'b1;
14558: pixelout<=1'b1;
14559: pixelout<=1'b1;
14560: pixelout<=1'b1;
14561: pixelout<=1'b1;
14562: pixelout<=1'b1;
14563: pixelout<=1'b1;
14564: pixelout<=1'b1;
14565: pixelout<=1'b1;
14566: pixelout<=1'b1;
14567: pixelout<=1'b1;
14568: pixelout<=1'b1;
14569: pixelout<=1'b1;
14570: pixelout<=1'b1;
14571: pixelout<=1'b1;
14572: pixelout<=1'b1;
14573: pixelout<=1'b1;
14574: pixelout<=1'b1;
14575: pixelout<=1'b1;
14576: pixelout<=1'b1;
14577: pixelout<=1'b1;
14578: pixelout<=1'b1;
14579: pixelout<=1'b1;
14580: pixelout<=1'b1;
14581: pixelout<=1'b1;
14582: pixelout<=1'b1;
14583: pixelout<=1'b1;
14584: pixelout<=1'b1;
14585: pixelout<=1'b1;
14586: pixelout<=1'b1;
14587: pixelout<=1'b1;
14588: pixelout<=1'b1;
14589: pixelout<=1'b1;
14590: pixelout<=1'b1;
14591: pixelout<=1'b1;
14592: pixelout<=1'b1;
14593: pixelout<=1'b1;
14594: pixelout<=1'b1;
14595: pixelout<=1'b1;
14596: pixelout<=1'b1;
14597: pixelout<=1'b1;
14598: pixelout<=1'b1;
14599: pixelout<=1'b1;
14600: pixelout<=1'b1;
14601: pixelout<=1'b1;
14602: pixelout<=1'b1;
14603: pixelout<=1'b1;
14604: pixelout<=1'b1;
14605: pixelout<=1'b1;
14606: pixelout<=1'b1;
14607: pixelout<=1'b0;
14608: pixelout<=1'b1;
14609: pixelout<=1'b1;
14610: pixelout<=1'b1;
14611: pixelout<=1'b1;
14612: pixelout<=1'b1;
14613: pixelout<=1'b1;
14614: pixelout<=1'b1;
14615: pixelout<=1'b1;
14616: pixelout<=1'b1;
14617: pixelout<=1'b1;
14618: pixelout<=1'b1;
14619: pixelout<=1'b1;
14620: pixelout<=1'b1;
14621: pixelout<=1'b1;
14622: pixelout<=1'b1;
14623: pixelout<=1'b1;
14624: pixelout<=1'b1;
14625: pixelout<=1'b1;
14626: pixelout<=1'b1;
14627: pixelout<=1'b1;
14628: pixelout<=1'b1;
14629: pixelout<=1'b1;
14630: pixelout<=1'b1;
14631: pixelout<=1'b1;
14632: pixelout<=1'b1;
14633: pixelout<=1'b1;
14634: pixelout<=1'b1;
14635: pixelout<=1'b1;
14636: pixelout<=1'b1;
14637: pixelout<=1'b1;
14638: pixelout<=1'b1;
14639: pixelout<=1'b1;
14640: pixelout<=1'b1;
14641: pixelout<=1'b1;
14642: pixelout<=1'b1;
14643: pixelout<=1'b1;
14644: pixelout<=1'b1;
14645: pixelout<=1'b1;
14646: pixelout<=1'b1;
14647: pixelout<=1'b1;
14648: pixelout<=1'b1;
14649: pixelout<=1'b1;
14650: pixelout<=1'b1;
14651: pixelout<=1'b1;
14652: pixelout<=1'b1;
14653: pixelout<=1'b1;
14654: pixelout<=1'b1;
14655: pixelout<=1'b1;
14656: pixelout<=1'b1;
14657: pixelout<=1'b1;
14658: pixelout<=1'b1;
14659: pixelout<=1'b1;
14660: pixelout<=1'b1;
14661: pixelout<=1'b1;
14662: pixelout<=1'b1;
14663: pixelout<=1'b1;
14664: pixelout<=1'b1;
14665: pixelout<=1'b1;
14666: pixelout<=1'b1;
14667: pixelout<=1'b1;
14668: pixelout<=1'b1;
14669: pixelout<=1'b1;
14670: pixelout<=1'b1;
14671: pixelout<=1'b1;
14672: pixelout<=1'b1;
14673: pixelout<=1'b1;
14674: pixelout<=1'b1;
14675: pixelout<=1'b1;
14676: pixelout<=1'b1;
14677: pixelout<=1'b1;
14678: pixelout<=1'b1;
14679: pixelout<=1'b1;
14680: pixelout<=1'b1;
14681: pixelout<=1'b1;
14682: pixelout<=1'b1;
14683: pixelout<=1'b1;
14684: pixelout<=1'b1;
14685: pixelout<=1'b1;
14686: pixelout<=1'b1;
14687: pixelout<=1'b1;
14688: pixelout<=1'b1;
14689: pixelout<=1'b1;
14690: pixelout<=1'b1;
14691: pixelout<=1'b1;
14692: pixelout<=1'b1;
14693: pixelout<=1'b1;
14694: pixelout<=1'b1;
14695: pixelout<=1'b1;
14696: pixelout<=1'b1;
14697: pixelout<=1'b1;
14698: pixelout<=1'b1;
14699: pixelout<=1'b1;
14700: pixelout<=1'b1;
14701: pixelout<=1'b1;
14702: pixelout<=1'b1;
14703: pixelout<=1'b1;
14704: pixelout<=1'b1;
14705: pixelout<=1'b1;
14706: pixelout<=1'b1;
14707: pixelout<=1'b1;
14708: pixelout<=1'b1;
14709: pixelout<=1'b1;
14710: pixelout<=1'b1;
14711: pixelout<=1'b1;
14712: pixelout<=1'b1;
14713: pixelout<=1'b1;
14714: pixelout<=1'b1;
14715: pixelout<=1'b1;
14716: pixelout<=1'b1;
14717: pixelout<=1'b1;
14718: pixelout<=1'b1;
14719: pixelout<=1'b1;
14720: pixelout<=1'b1;
14721: pixelout<=1'b1;
14722: pixelout<=1'b1;
14723: pixelout<=1'b1;
14724: pixelout<=1'b1;
14725: pixelout<=1'b1;
14726: pixelout<=1'b1;
14727: pixelout<=1'b1;
14728: pixelout<=1'b1;
14729: pixelout<=1'b1;
14730: pixelout<=1'b1;
14731: pixelout<=1'b1;
14732: pixelout<=1'b1;
14733: pixelout<=1'b1;
14734: pixelout<=1'b1;
14735: pixelout<=1'b1;
14736: pixelout<=1'b1;
14737: pixelout<=1'b1;
14738: pixelout<=1'b1;
14739: pixelout<=1'b1;
14740: pixelout<=1'b1;
14741: pixelout<=1'b1;
14742: pixelout<=1'b1;
14743: pixelout<=1'b1;
14744: pixelout<=1'b1;
14745: pixelout<=1'b1;
14746: pixelout<=1'b1;
14747: pixelout<=1'b1;
14748: pixelout<=1'b1;
14749: pixelout<=1'b1;
14750: pixelout<=1'b1;
14751: pixelout<=1'b1;
14752: pixelout<=1'b1;
14753: pixelout<=1'b1;
14754: pixelout<=1'b1;
14755: pixelout<=1'b1;
14756: pixelout<=1'b1;
14757: pixelout<=1'b1;
14758: pixelout<=1'b1;
14759: pixelout<=1'b1;
14760: pixelout<=1'b1;
14761: pixelout<=1'b1;
14762: pixelout<=1'b1;
14763: pixelout<=1'b1;
14764: pixelout<=1'b1;
14765: pixelout<=1'b1;
14766: pixelout<=1'b1;
14767: pixelout<=1'b1;
14768: pixelout<=1'b1;
14769: pixelout<=1'b1;
14770: pixelout<=1'b1;
14771: pixelout<=1'b1;
14772: pixelout<=1'b1;
14773: pixelout<=1'b1;
14774: pixelout<=1'b1;
14775: pixelout<=1'b1;
14776: pixelout<=1'b1;
14777: pixelout<=1'b1;
14778: pixelout<=1'b1;
14779: pixelout<=1'b1;
14780: pixelout<=1'b1;
14781: pixelout<=1'b1;
14782: pixelout<=1'b1;
14783: pixelout<=1'b1;
14784: pixelout<=1'b1;
14785: pixelout<=1'b1;
14786: pixelout<=1'b1;
14787: pixelout<=1'b1;
14788: pixelout<=1'b1;
14789: pixelout<=1'b1;
14790: pixelout<=1'b1;
14791: pixelout<=1'b1;
14792: pixelout<=1'b1;
14793: pixelout<=1'b1;
14794: pixelout<=1'b1;
14795: pixelout<=1'b1;
14796: pixelout<=1'b1;
14797: pixelout<=1'b1;
14798: pixelout<=1'b1;
14799: pixelout<=1'b1;
14800: pixelout<=1'b1;
14801: pixelout<=1'b1;
14802: pixelout<=1'b1;
14803: pixelout<=1'b1;
14804: pixelout<=1'b1;
14805: pixelout<=1'b1;
14806: pixelout<=1'b1;
14807: pixelout<=1'b1;
14808: pixelout<=1'b1;
14809: pixelout<=1'b1;
14810: pixelout<=1'b1;
14811: pixelout<=1'b1;
14812: pixelout<=1'b1;
14813: pixelout<=1'b1;
14814: pixelout<=1'b1;
14815: pixelout<=1'b1;
14816: pixelout<=1'b1;
14817: pixelout<=1'b1;
14818: pixelout<=1'b1;
14819: pixelout<=1'b1;
14820: pixelout<=1'b1;
14821: pixelout<=1'b1;
14822: pixelout<=1'b1;
14823: pixelout<=1'b1;
14824: pixelout<=1'b1;
14825: pixelout<=1'b1;
14826: pixelout<=1'b1;
14827: pixelout<=1'b1;
14828: pixelout<=1'b1;
14829: pixelout<=1'b1;
14830: pixelout<=1'b1;
14831: pixelout<=1'b1;
14832: pixelout<=1'b1;
14833: pixelout<=1'b1;
14834: pixelout<=1'b1;
14835: pixelout<=1'b1;
14836: pixelout<=1'b1;
14837: pixelout<=1'b1;
14838: pixelout<=1'b1;
14839: pixelout<=1'b1;
14840: pixelout<=1'b1;
14841: pixelout<=1'b1;
14842: pixelout<=1'b1;
14843: pixelout<=1'b1;
14844: pixelout<=1'b1;
14845: pixelout<=1'b1;
14846: pixelout<=1'b1;
14847: pixelout<=1'b1;
14848: pixelout<=1'b1;
14849: pixelout<=1'b1;
14850: pixelout<=1'b1;
14851: pixelout<=1'b1;
14852: pixelout<=1'b1;
14853: pixelout<=1'b1;
14854: pixelout<=1'b1;
14855: pixelout<=1'b1;
14856: pixelout<=1'b1;
14857: pixelout<=1'b1;
14858: pixelout<=1'b1;
14859: pixelout<=1'b1;
14860: pixelout<=1'b1;
14861: pixelout<=1'b1;
14862: pixelout<=1'b1;
14863: pixelout<=1'b1;
14864: pixelout<=1'b1;
14865: pixelout<=1'b1;
14866: pixelout<=1'b1;
14867: pixelout<=1'b1;
14868: pixelout<=1'b1;
14869: pixelout<=1'b1;
14870: pixelout<=1'b1;
14871: pixelout<=1'b1;
14872: pixelout<=1'b1;
14873: pixelout<=1'b1;
14874: pixelout<=1'b1;
14875: pixelout<=1'b1;
14876: pixelout<=1'b1;
14877: pixelout<=1'b1;
14878: pixelout<=1'b1;
14879: pixelout<=1'b1;
14880: pixelout<=1'b1;
14881: pixelout<=1'b1;
14882: pixelout<=1'b1;
14883: pixelout<=1'b1;
14884: pixelout<=1'b1;
14885: pixelout<=1'b1;
14886: pixelout<=1'b1;
14887: pixelout<=1'b1;
14888: pixelout<=1'b1;
14889: pixelout<=1'b1;
14890: pixelout<=1'b1;
14891: pixelout<=1'b1;
14892: pixelout<=1'b1;
14893: pixelout<=1'b1;
14894: pixelout<=1'b1;
14895: pixelout<=1'b1;
14896: pixelout<=1'b1;
14897: pixelout<=1'b1;
14898: pixelout<=1'b1;
14899: pixelout<=1'b1;
14900: pixelout<=1'b1;
14901: pixelout<=1'b1;
14902: pixelout<=1'b1;
14903: pixelout<=1'b1;
14904: pixelout<=1'b1;
14905: pixelout<=1'b1;
14906: pixelout<=1'b1;
14907: pixelout<=1'b1;
14908: pixelout<=1'b1;
14909: pixelout<=1'b1;
14910: pixelout<=1'b1;
14911: pixelout<=1'b1;
14912: pixelout<=1'b1;
14913: pixelout<=1'b1;
14914: pixelout<=1'b1;
14915: pixelout<=1'b1;
14916: pixelout<=1'b1;
14917: pixelout<=1'b1;
14918: pixelout<=1'b1;
14919: pixelout<=1'b1;
14920: pixelout<=1'b1;
14921: pixelout<=1'b1;
14922: pixelout<=1'b1;
14923: pixelout<=1'b1;
14924: pixelout<=1'b1;
14925: pixelout<=1'b1;
14926: pixelout<=1'b1;
14927: pixelout<=1'b1;
14928: pixelout<=1'b1;
14929: pixelout<=1'b1;
14930: pixelout<=1'b1;
14931: pixelout<=1'b1;
14932: pixelout<=1'b1;
14933: pixelout<=1'b1;
14934: pixelout<=1'b1;
14935: pixelout<=1'b1;
14936: pixelout<=1'b1;
14937: pixelout<=1'b1;
14938: pixelout<=1'b1;
14939: pixelout<=1'b1;
14940: pixelout<=1'b1;
14941: pixelout<=1'b1;
14942: pixelout<=1'b1;
14943: pixelout<=1'b1;
14944: pixelout<=1'b1;
14945: pixelout<=1'b1;
14946: pixelout<=1'b1;
14947: pixelout<=1'b1;
14948: pixelout<=1'b1;
14949: pixelout<=1'b1;
14950: pixelout<=1'b1;
14951: pixelout<=1'b1;
14952: pixelout<=1'b1;
14953: pixelout<=1'b1;
14954: pixelout<=1'b1;
14955: pixelout<=1'b1;
14956: pixelout<=1'b1;
14957: pixelout<=1'b1;
14958: pixelout<=1'b1;
14959: pixelout<=1'b1;
14960: pixelout<=1'b1;
14961: pixelout<=1'b1;
14962: pixelout<=1'b1;
14963: pixelout<=1'b1;
14964: pixelout<=1'b1;
14965: pixelout<=1'b1;
14966: pixelout<=1'b1;
14967: pixelout<=1'b1;
14968: pixelout<=1'b1;
14969: pixelout<=1'b1;
14970: pixelout<=1'b1;
14971: pixelout<=1'b1;
14972: pixelout<=1'b1;
14973: pixelout<=1'b1;
14974: pixelout<=1'b1;
14975: pixelout<=1'b1;
14976: pixelout<=1'b1;
14977: pixelout<=1'b1;
14978: pixelout<=1'b1;
14979: pixelout<=1'b1;
14980: pixelout<=1'b1;
14981: pixelout<=1'b1;
14982: pixelout<=1'b1;
14983: pixelout<=1'b1;
14984: pixelout<=1'b1;
14985: pixelout<=1'b1;
14986: pixelout<=1'b1;
14987: pixelout<=1'b1;
14988: pixelout<=1'b1;
14989: pixelout<=1'b1;
14990: pixelout<=1'b1;
14991: pixelout<=1'b1;
14992: pixelout<=1'b1;
14993: pixelout<=1'b1;
14994: pixelout<=1'b1;
14995: pixelout<=1'b1;
14996: pixelout<=1'b1;
14997: pixelout<=1'b1;
14998: pixelout<=1'b1;
14999: pixelout<=1'b1;
15000: pixelout<=1'b1;
15001: pixelout<=1'b1;
15002: pixelout<=1'b1;
15003: pixelout<=1'b1;
15004: pixelout<=1'b1;
15005: pixelout<=1'b1;
15006: pixelout<=1'b1;
15007: pixelout<=1'b1;
15008: pixelout<=1'b1;
15009: pixelout<=1'b1;
15010: pixelout<=1'b1;
15011: pixelout<=1'b1;
15012: pixelout<=1'b1;
15013: pixelout<=1'b1;
15014: pixelout<=1'b1;
15015: pixelout<=1'b1;
15016: pixelout<=1'b1;
15017: pixelout<=1'b1;
15018: pixelout<=1'b1;
15019: pixelout<=1'b1;
15020: pixelout<=1'b1;
15021: pixelout<=1'b1;
15022: pixelout<=1'b1;
15023: pixelout<=1'b1;
15024: pixelout<=1'b1;
15025: pixelout<=1'b1;
15026: pixelout<=1'b1;
15027: pixelout<=1'b1;
15028: pixelout<=1'b1;
15029: pixelout<=1'b1;
15030: pixelout<=1'b1;
15031: pixelout<=1'b1;
15032: pixelout<=1'b1;
15033: pixelout<=1'b1;
15034: pixelout<=1'b1;
15035: pixelout<=1'b1;
15036: pixelout<=1'b1;
15037: pixelout<=1'b1;
15038: pixelout<=1'b1;
15039: pixelout<=1'b1;
15040: pixelout<=1'b1;
15041: pixelout<=1'b1;
15042: pixelout<=1'b1;
15043: pixelout<=1'b1;
15044: pixelout<=1'b1;
15045: pixelout<=1'b1;
15046: pixelout<=1'b1;
15047: pixelout<=1'b1;
15048: pixelout<=1'b1;
15049: pixelout<=1'b1;
15050: pixelout<=1'b1;
15051: pixelout<=1'b1;
15052: pixelout<=1'b1;
15053: pixelout<=1'b1;
15054: pixelout<=1'b1;
15055: pixelout<=1'b1;
15056: pixelout<=1'b1;
15057: pixelout<=1'b1;
15058: pixelout<=1'b1;
15059: pixelout<=1'b1;
15060: pixelout<=1'b1;
15061: pixelout<=1'b1;
15062: pixelout<=1'b1;
15063: pixelout<=1'b1;
15064: pixelout<=1'b1;
15065: pixelout<=1'b1;
15066: pixelout<=1'b1;
15067: pixelout<=1'b1;
15068: pixelout<=1'b1;
15069: pixelout<=1'b1;
15070: pixelout<=1'b1;
15071: pixelout<=1'b1;
15072: pixelout<=1'b1;
15073: pixelout<=1'b1;
15074: pixelout<=1'b1;
15075: pixelout<=1'b1;
15076: pixelout<=1'b1;
15077: pixelout<=1'b1;
15078: pixelout<=1'b1;
15079: pixelout<=1'b1;
15080: pixelout<=1'b1;
15081: pixelout<=1'b1;
15082: pixelout<=1'b1;
15083: pixelout<=1'b1;
15084: pixelout<=1'b1;
15085: pixelout<=1'b1;
15086: pixelout<=1'b1;
15087: pixelout<=1'b1;
15088: pixelout<=1'b1;
15089: pixelout<=1'b1;
15090: pixelout<=1'b1;
15091: pixelout<=1'b1;
15092: pixelout<=1'b1;
15093: pixelout<=1'b1;
15094: pixelout<=1'b1;
15095: pixelout<=1'b1;
15096: pixelout<=1'b1;
15097: pixelout<=1'b1;
15098: pixelout<=1'b1;
15099: pixelout<=1'b1;
15100: pixelout<=1'b1;
15101: pixelout<=1'b1;
15102: pixelout<=1'b1;
15103: pixelout<=1'b1;
15104: pixelout<=1'b1;
15105: pixelout<=1'b1;
15106: pixelout<=1'b1;
15107: pixelout<=1'b1;
15108: pixelout<=1'b1;
15109: pixelout<=1'b1;
15110: pixelout<=1'b1;
15111: pixelout<=1'b1;
15112: pixelout<=1'b1;
15113: pixelout<=1'b1;
15114: pixelout<=1'b1;
15115: pixelout<=1'b1;
15116: pixelout<=1'b1;
15117: pixelout<=1'b1;
15118: pixelout<=1'b1;
15119: pixelout<=1'b1;
15120: pixelout<=1'b1;
15121: pixelout<=1'b1;
15122: pixelout<=1'b1;
15123: pixelout<=1'b1;
15124: pixelout<=1'b1;
15125: pixelout<=1'b1;
15126: pixelout<=1'b1;
15127: pixelout<=1'b1;
15128: pixelout<=1'b1;
15129: pixelout<=1'b1;
15130: pixelout<=1'b1;
15131: pixelout<=1'b1;
15132: pixelout<=1'b1;
15133: pixelout<=1'b1;
15134: pixelout<=1'b1;
15135: pixelout<=1'b1;
15136: pixelout<=1'b1;
15137: pixelout<=1'b1;
15138: pixelout<=1'b1;
15139: pixelout<=1'b1;
15140: pixelout<=1'b1;
15141: pixelout<=1'b1;
15142: pixelout<=1'b1;
15143: pixelout<=1'b1;
15144: pixelout<=1'b1;
15145: pixelout<=1'b1;
15146: pixelout<=1'b1;
15147: pixelout<=1'b1;
15148: pixelout<=1'b1;
15149: pixelout<=1'b1;
15150: pixelout<=1'b1;
15151: pixelout<=1'b1;
15152: pixelout<=1'b1;
15153: pixelout<=1'b1;
15154: pixelout<=1'b1;
15155: pixelout<=1'b1;
15156: pixelout<=1'b1;
15157: pixelout<=1'b1;
15158: pixelout<=1'b1;
15159: pixelout<=1'b1;
15160: pixelout<=1'b1;
15161: pixelout<=1'b1;
15162: pixelout<=1'b1;
15163: pixelout<=1'b1;
15164: pixelout<=1'b1;
15165: pixelout<=1'b1;
15166: pixelout<=1'b1;
15167: pixelout<=1'b1;
15168: pixelout<=1'b1;
15169: pixelout<=1'b1;
15170: pixelout<=1'b1;
15171: pixelout<=1'b1;
15172: pixelout<=1'b1;
15173: pixelout<=1'b1;
15174: pixelout<=1'b1;
15175: pixelout<=1'b1;
15176: pixelout<=1'b1;
15177: pixelout<=1'b1;
15178: pixelout<=1'b1;
15179: pixelout<=1'b1;
15180: pixelout<=1'b1;
15181: pixelout<=1'b1;
15182: pixelout<=1'b1;
15183: pixelout<=1'b1;
15184: pixelout<=1'b1;
15185: pixelout<=1'b1;
15186: pixelout<=1'b1;
15187: pixelout<=1'b1;
15188: pixelout<=1'b1;
15189: pixelout<=1'b1;
15190: pixelout<=1'b1;
15191: pixelout<=1'b1;
15192: pixelout<=1'b1;
15193: pixelout<=1'b1;
15194: pixelout<=1'b1;
15195: pixelout<=1'b1;
15196: pixelout<=1'b1;
15197: pixelout<=1'b1;
15198: pixelout<=1'b1;
15199: pixelout<=1'b1;
15200: pixelout<=1'b1;
15201: pixelout<=1'b1;
15202: pixelout<=1'b1;
15203: pixelout<=1'b1;
15204: pixelout<=1'b1;
15205: pixelout<=1'b1;
15206: pixelout<=1'b1;
15207: pixelout<=1'b1;
15208: pixelout<=1'b1;
15209: pixelout<=1'b1;
15210: pixelout<=1'b1;
15211: pixelout<=1'b1;
15212: pixelout<=1'b1;
15213: pixelout<=1'b1;
15214: pixelout<=1'b1;
15215: pixelout<=1'b1;
15216: pixelout<=1'b1;
15217: pixelout<=1'b1;
15218: pixelout<=1'b1;
15219: pixelout<=1'b1;
15220: pixelout<=1'b1;
15221: pixelout<=1'b1;
15222: pixelout<=1'b1;
15223: pixelout<=1'b1;
15224: pixelout<=1'b1;
15225: pixelout<=1'b1;
15226: pixelout<=1'b1;
15227: pixelout<=1'b1;
15228: pixelout<=1'b1;
15229: pixelout<=1'b1;
15230: pixelout<=1'b1;
15231: pixelout<=1'b1;
15232: pixelout<=1'b1;
15233: pixelout<=1'b1;
15234: pixelout<=1'b1;
15235: pixelout<=1'b1;
15236: pixelout<=1'b1;
15237: pixelout<=1'b1;
15238: pixelout<=1'b1;
15239: pixelout<=1'b1;
15240: pixelout<=1'b1;
15241: pixelout<=1'b1;
15242: pixelout<=1'b1;
15243: pixelout<=1'b1;
15244: pixelout<=1'b1;
15245: pixelout<=1'b1;
15246: pixelout<=1'b1;
15247: pixelout<=1'b1;
15248: pixelout<=1'b1;
15249: pixelout<=1'b1;
15250: pixelout<=1'b1;
15251: pixelout<=1'b1;
15252: pixelout<=1'b1;
15253: pixelout<=1'b1;
15254: pixelout<=1'b1;
15255: pixelout<=1'b1;
15256: pixelout<=1'b1;
15257: pixelout<=1'b1;
15258: pixelout<=1'b1;
15259: pixelout<=1'b1;
15260: pixelout<=1'b1;
15261: pixelout<=1'b1;
15262: pixelout<=1'b1;
15263: pixelout<=1'b1;
15264: pixelout<=1'b1;
15265: pixelout<=1'b1;
15266: pixelout<=1'b1;
15267: pixelout<=1'b1;
15268: pixelout<=1'b1;
15269: pixelout<=1'b1;
15270: pixelout<=1'b1;
15271: pixelout<=1'b1;
15272: pixelout<=1'b1;
15273: pixelout<=1'b1;
15274: pixelout<=1'b1;
15275: pixelout<=1'b1;
15276: pixelout<=1'b1;
15277: pixelout<=1'b1;
15278: pixelout<=1'b1;
15279: pixelout<=1'b1;
15280: pixelout<=1'b1;
15281: pixelout<=1'b1;
15282: pixelout<=1'b1;
15283: pixelout<=1'b1;
15284: pixelout<=1'b1;
15285: pixelout<=1'b1;
15286: pixelout<=1'b1;
15287: pixelout<=1'b1;
15288: pixelout<=1'b1;
15289: pixelout<=1'b1;
15290: pixelout<=1'b1;
15291: pixelout<=1'b1;
15292: pixelout<=1'b1;
15293: pixelout<=1'b1;
15294: pixelout<=1'b1;
15295: pixelout<=1'b1;
15296: pixelout<=1'b1;
15297: pixelout<=1'b1;
15298: pixelout<=1'b1;
15299: pixelout<=1'b1;
15300: pixelout<=1'b1;
15301: pixelout<=1'b1;
15302: pixelout<=1'b1;
15303: pixelout<=1'b1;
15304: pixelout<=1'b1;
15305: pixelout<=1'b1;
15306: pixelout<=1'b1;
15307: pixelout<=1'b1;
15308: pixelout<=1'b1;
15309: pixelout<=1'b1;
15310: pixelout<=1'b1;
15311: pixelout<=1'b1;
15312: pixelout<=1'b1;
15313: pixelout<=1'b1;
15314: pixelout<=1'b1;
15315: pixelout<=1'b1;
15316: pixelout<=1'b1;
15317: pixelout<=1'b1;
15318: pixelout<=1'b1;
15319: pixelout<=1'b1;
15320: pixelout<=1'b1;
15321: pixelout<=1'b1;
15322: pixelout<=1'b1;
15323: pixelout<=1'b1;
15324: pixelout<=1'b1;
15325: pixelout<=1'b1;
15326: pixelout<=1'b1;
15327: pixelout<=1'b1;
15328: pixelout<=1'b1;
15329: pixelout<=1'b1;
15330: pixelout<=1'b1;
15331: pixelout<=1'b1;
15332: pixelout<=1'b1;
15333: pixelout<=1'b1;
15334: pixelout<=1'b1;
15335: pixelout<=1'b1;
15336: pixelout<=1'b1;
15337: pixelout<=1'b1;
15338: pixelout<=1'b1;
15339: pixelout<=1'b1;
15340: pixelout<=1'b1;
15341: pixelout<=1'b1;
15342: pixelout<=1'b1;
15343: pixelout<=1'b1;
15344: pixelout<=1'b1;
15345: pixelout<=1'b1;
15346: pixelout<=1'b1;
15347: pixelout<=1'b1;
15348: pixelout<=1'b1;
15349: pixelout<=1'b1;
15350: pixelout<=1'b1;
15351: pixelout<=1'b1;
15352: pixelout<=1'b1;
15353: pixelout<=1'b1;
15354: pixelout<=1'b1;
15355: pixelout<=1'b1;
15356: pixelout<=1'b1;
15357: pixelout<=1'b1;
15358: pixelout<=1'b1;
15359: pixelout<=1'b1;
15360: pixelout<=1'b1;
15361: pixelout<=1'b1;
15362: pixelout<=1'b1;
15363: pixelout<=1'b1;
15364: pixelout<=1'b1;
15365: pixelout<=1'b1;
15366: pixelout<=1'b1;
15367: pixelout<=1'b1;
15368: pixelout<=1'b1;
15369: pixelout<=1'b1;
15370: pixelout<=1'b1;
15371: pixelout<=1'b1;
15372: pixelout<=1'b1;
15373: pixelout<=1'b1;
15374: pixelout<=1'b1;
15375: pixelout<=1'b1;
15376: pixelout<=1'b1;
15377: pixelout<=1'b1;
15378: pixelout<=1'b1;
15379: pixelout<=1'b1;
15380: pixelout<=1'b1;
15381: pixelout<=1'b1;
15382: pixelout<=1'b1;
15383: pixelout<=1'b1;
15384: pixelout<=1'b1;
15385: pixelout<=1'b1;
15386: pixelout<=1'b1;
15387: pixelout<=1'b1;
15388: pixelout<=1'b1;
15389: pixelout<=1'b1;
15390: pixelout<=1'b1;
15391: pixelout<=1'b1;
15392: pixelout<=1'b1;
15393: pixelout<=1'b1;
15394: pixelout<=1'b1;
15395: pixelout<=1'b1;
15396: pixelout<=1'b1;
15397: pixelout<=1'b1;
15398: pixelout<=1'b1;
15399: pixelout<=1'b1;
15400: pixelout<=1'b1;
15401: pixelout<=1'b1;
15402: pixelout<=1'b1;
15403: pixelout<=1'b1;
15404: pixelout<=1'b1;
15405: pixelout<=1'b1;
15406: pixelout<=1'b1;
15407: pixelout<=1'b1;
15408: pixelout<=1'b1;
15409: pixelout<=1'b1;
15410: pixelout<=1'b1;
15411: pixelout<=1'b1;
15412: pixelout<=1'b1;
15413: pixelout<=1'b1;
15414: pixelout<=1'b1;
15415: pixelout<=1'b1;
15416: pixelout<=1'b1;
15417: pixelout<=1'b1;
15418: pixelout<=1'b1;
15419: pixelout<=1'b1;
15420: pixelout<=1'b1;
15421: pixelout<=1'b1;
15422: pixelout<=1'b1;
15423: pixelout<=1'b1;
15424: pixelout<=1'b1;
15425: pixelout<=1'b1;
15426: pixelout<=1'b1;
15427: pixelout<=1'b1;
15428: pixelout<=1'b1;
15429: pixelout<=1'b1;
15430: pixelout<=1'b1;
15431: pixelout<=1'b1;
15432: pixelout<=1'b1;
15433: pixelout<=1'b1;
15434: pixelout<=1'b1;
15435: pixelout<=1'b1;
15436: pixelout<=1'b1;
15437: pixelout<=1'b1;
15438: pixelout<=1'b1;
15439: pixelout<=1'b1;
15440: pixelout<=1'b1;
15441: pixelout<=1'b1;
15442: pixelout<=1'b1;
15443: pixelout<=1'b1;
15444: pixelout<=1'b1;
15445: pixelout<=1'b1;
15446: pixelout<=1'b1;
15447: pixelout<=1'b1;
15448: pixelout<=1'b1;
15449: pixelout<=1'b1;
15450: pixelout<=1'b1;
15451: pixelout<=1'b1;
15452: pixelout<=1'b1;
15453: pixelout<=1'b1;
15454: pixelout<=1'b1;
15455: pixelout<=1'b1;
15456: pixelout<=1'b1;
15457: pixelout<=1'b1;
15458: pixelout<=1'b1;
15459: pixelout<=1'b1;
15460: pixelout<=1'b1;
15461: pixelout<=1'b1;
15462: pixelout<=1'b1;
15463: pixelout<=1'b1;
15464: pixelout<=1'b1;
15465: pixelout<=1'b1;
15466: pixelout<=1'b1;
15467: pixelout<=1'b1;
15468: pixelout<=1'b1;
15469: pixelout<=1'b1;
15470: pixelout<=1'b1;
15471: pixelout<=1'b1;
15472: pixelout<=1'b1;
15473: pixelout<=1'b1;
15474: pixelout<=1'b1;
15475: pixelout<=1'b1;
15476: pixelout<=1'b1;
15477: pixelout<=1'b1;
15478: pixelout<=1'b1;
15479: pixelout<=1'b1;
15480: pixelout<=1'b1;
15481: pixelout<=1'b1;
15482: pixelout<=1'b1;
15483: pixelout<=1'b1;
15484: pixelout<=1'b1;
15485: pixelout<=1'b1;
15486: pixelout<=1'b1;
15487: pixelout<=1'b1;
15488: pixelout<=1'b1;
15489: pixelout<=1'b1;
15490: pixelout<=1'b1;
15491: pixelout<=1'b1;
15492: pixelout<=1'b1;
15493: pixelout<=1'b1;
15494: pixelout<=1'b1;
15495: pixelout<=1'b1;
15496: pixelout<=1'b1;
15497: pixelout<=1'b1;
15498: pixelout<=1'b1;
15499: pixelout<=1'b1;
15500: pixelout<=1'b1;
15501: pixelout<=1'b1;
15502: pixelout<=1'b1;
15503: pixelout<=1'b1;
15504: pixelout<=1'b1;
15505: pixelout<=1'b1;
15506: pixelout<=1'b1;
15507: pixelout<=1'b1;
15508: pixelout<=1'b1;
15509: pixelout<=1'b1;
15510: pixelout<=1'b1;
15511: pixelout<=1'b1;
15512: pixelout<=1'b1;
15513: pixelout<=1'b1;
15514: pixelout<=1'b1;
15515: pixelout<=1'b1;
15516: pixelout<=1'b1;
15517: pixelout<=1'b1;
15518: pixelout<=1'b1;
15519: pixelout<=1'b1;
15520: pixelout<=1'b1;
15521: pixelout<=1'b1;
15522: pixelout<=1'b1;
15523: pixelout<=1'b1;
15524: pixelout<=1'b1;
15525: pixelout<=1'b1;
15526: pixelout<=1'b1;
15527: pixelout<=1'b1;
15528: pixelout<=1'b1;
15529: pixelout<=1'b1;
15530: pixelout<=1'b1;
15531: pixelout<=1'b1;
15532: pixelout<=1'b1;
15533: pixelout<=1'b1;
15534: pixelout<=1'b1;
15535: pixelout<=1'b1;
15536: pixelout<=1'b1;
15537: pixelout<=1'b1;
15538: pixelout<=1'b1;
15539: pixelout<=1'b1;
15540: pixelout<=1'b1;
15541: pixelout<=1'b1;
15542: pixelout<=1'b1;
15543: pixelout<=1'b1;
15544: pixelout<=1'b1;
15545: pixelout<=1'b1;
15546: pixelout<=1'b1;
15547: pixelout<=1'b1;
15548: pixelout<=1'b1;
15549: pixelout<=1'b1;
15550: pixelout<=1'b1;
15551: pixelout<=1'b1;
15552: pixelout<=1'b1;
15553: pixelout<=1'b1;
15554: pixelout<=1'b1;
15555: pixelout<=1'b1;
15556: pixelout<=1'b1;
15557: pixelout<=1'b1;
15558: pixelout<=1'b1;
15559: pixelout<=1'b1;
15560: pixelout<=1'b1;
15561: pixelout<=1'b1;
15562: pixelout<=1'b1;
15563: pixelout<=1'b1;
15564: pixelout<=1'b1;
15565: pixelout<=1'b1;
15566: pixelout<=1'b1;
15567: pixelout<=1'b1;
15568: pixelout<=1'b1;
15569: pixelout<=1'b1;
15570: pixelout<=1'b1;
15571: pixelout<=1'b1;
15572: pixelout<=1'b1;
15573: pixelout<=1'b1;
15574: pixelout<=1'b1;
15575: pixelout<=1'b1;
15576: pixelout<=1'b1;
15577: pixelout<=1'b1;
15578: pixelout<=1'b1;
15579: pixelout<=1'b1;
15580: pixelout<=1'b1;
15581: pixelout<=1'b1;
15582: pixelout<=1'b1;
15583: pixelout<=1'b1;
15584: pixelout<=1'b1;
15585: pixelout<=1'b1;
15586: pixelout<=1'b1;
15587: pixelout<=1'b1;
15588: pixelout<=1'b1;
15589: pixelout<=1'b1;
15590: pixelout<=1'b1;
15591: pixelout<=1'b1;
15592: pixelout<=1'b1;
15593: pixelout<=1'b1;
15594: pixelout<=1'b1;
15595: pixelout<=1'b1;
15596: pixelout<=1'b1;
15597: pixelout<=1'b1;
15598: pixelout<=1'b1;
15599: pixelout<=1'b1;
15600: pixelout<=1'b1;
15601: pixelout<=1'b1;
15602: pixelout<=1'b1;
15603: pixelout<=1'b1;
15604: pixelout<=1'b1;
15605: pixelout<=1'b1;
15606: pixelout<=1'b1;
15607: pixelout<=1'b1;
15608: pixelout<=1'b1;
15609: pixelout<=1'b1;
15610: pixelout<=1'b1;
15611: pixelout<=1'b1;
15612: pixelout<=1'b1;
15613: pixelout<=1'b1;
15614: pixelout<=1'b1;
15615: pixelout<=1'b1;
15616: pixelout<=1'b1;
15617: pixelout<=1'b1;
15618: pixelout<=1'b1;
15619: pixelout<=1'b1;
15620: pixelout<=1'b1;
15621: pixelout<=1'b1;
15622: pixelout<=1'b1;
15623: pixelout<=1'b1;
15624: pixelout<=1'b1;
15625: pixelout<=1'b1;
15626: pixelout<=1'b1;
15627: pixelout<=1'b1;
15628: pixelout<=1'b1;
15629: pixelout<=1'b1;
15630: pixelout<=1'b1;
15631: pixelout<=1'b1;
15632: pixelout<=1'b1;
15633: pixelout<=1'b1;
15634: pixelout<=1'b1;
15635: pixelout<=1'b1;
15636: pixelout<=1'b1;
15637: pixelout<=1'b1;
15638: pixelout<=1'b1;
15639: pixelout<=1'b1;
15640: pixelout<=1'b1;
15641: pixelout<=1'b1;
15642: pixelout<=1'b1;
15643: pixelout<=1'b1;
15644: pixelout<=1'b1;
15645: pixelout<=1'b1;
15646: pixelout<=1'b1;
15647: pixelout<=1'b1;
15648: pixelout<=1'b1;
15649: pixelout<=1'b1;
15650: pixelout<=1'b1;
15651: pixelout<=1'b1;
15652: pixelout<=1'b1;
15653: pixelout<=1'b1;
15654: pixelout<=1'b1;
15655: pixelout<=1'b1;
15656: pixelout<=1'b1;
15657: pixelout<=1'b1;
15658: pixelout<=1'b1;
15659: pixelout<=1'b1;
15660: pixelout<=1'b1;
15661: pixelout<=1'b1;
15662: pixelout<=1'b1;
15663: pixelout<=1'b1;
15664: pixelout<=1'b1;
15665: pixelout<=1'b1;
15666: pixelout<=1'b1;
15667: pixelout<=1'b1;
15668: pixelout<=1'b1;
15669: pixelout<=1'b1;
15670: pixelout<=1'b1;
15671: pixelout<=1'b1;
15672: pixelout<=1'b1;
15673: pixelout<=1'b1;
15674: pixelout<=1'b1;
15675: pixelout<=1'b1;
15676: pixelout<=1'b1;
15677: pixelout<=1'b1;
15678: pixelout<=1'b1;
15679: pixelout<=1'b1;
15680: pixelout<=1'b1;
15681: pixelout<=1'b1;
15682: pixelout<=1'b1;
15683: pixelout<=1'b1;
15684: pixelout<=1'b1;
15685: pixelout<=1'b1;
15686: pixelout<=1'b1;
15687: pixelout<=1'b1;
15688: pixelout<=1'b1;
15689: pixelout<=1'b1;
15690: pixelout<=1'b1;
15691: pixelout<=1'b1;
15692: pixelout<=1'b1;
15693: pixelout<=1'b1;
15694: pixelout<=1'b1;
15695: pixelout<=1'b1;
15696: pixelout<=1'b1;
15697: pixelout<=1'b1;
15698: pixelout<=1'b1;
15699: pixelout<=1'b1;
15700: pixelout<=1'b1;
15701: pixelout<=1'b1;
15702: pixelout<=1'b1;
15703: pixelout<=1'b1;
15704: pixelout<=1'b1;
15705: pixelout<=1'b1;
15706: pixelout<=1'b1;
15707: pixelout<=1'b1;
15708: pixelout<=1'b1;
15709: pixelout<=1'b1;
15710: pixelout<=1'b1;
15711: pixelout<=1'b1;
15712: pixelout<=1'b1;
15713: pixelout<=1'b1;
15714: pixelout<=1'b1;
15715: pixelout<=1'b1;
15716: pixelout<=1'b1;
15717: pixelout<=1'b1;
15718: pixelout<=1'b1;
15719: pixelout<=1'b1;
15720: pixelout<=1'b1;
15721: pixelout<=1'b1;
15722: pixelout<=1'b1;
15723: pixelout<=1'b1;
15724: pixelout<=1'b1;
15725: pixelout<=1'b1;
15726: pixelout<=1'b1;
15727: pixelout<=1'b1;
15728: pixelout<=1'b1;
15729: pixelout<=1'b1;
15730: pixelout<=1'b1;
15731: pixelout<=1'b1;
15732: pixelout<=1'b1;
15733: pixelout<=1'b1;
15734: pixelout<=1'b1;
15735: pixelout<=1'b1;
15736: pixelout<=1'b1;
15737: pixelout<=1'b1;
15738: pixelout<=1'b1;
15739: pixelout<=1'b1;
15740: pixelout<=1'b1;
15741: pixelout<=1'b1;
15742: pixelout<=1'b1;
15743: pixelout<=1'b1;
15744: pixelout<=1'b1;
15745: pixelout<=1'b1;
15746: pixelout<=1'b1;
15747: pixelout<=1'b1;
15748: pixelout<=1'b1;
15749: pixelout<=1'b1;
15750: pixelout<=1'b1;
15751: pixelout<=1'b1;
15752: pixelout<=1'b1;
15753: pixelout<=1'b1;
15754: pixelout<=1'b1;
15755: pixelout<=1'b1;
15756: pixelout<=1'b1;
15757: pixelout<=1'b1;
15758: pixelout<=1'b1;
15759: pixelout<=1'b1;
15760: pixelout<=1'b1;
15761: pixelout<=1'b1;
15762: pixelout<=1'b1;
15763: pixelout<=1'b1;
15764: pixelout<=1'b1;
15765: pixelout<=1'b1;
15766: pixelout<=1'b1;
15767: pixelout<=1'b1;
15768: pixelout<=1'b1;
15769: pixelout<=1'b1;
15770: pixelout<=1'b1;
15771: pixelout<=1'b1;
15772: pixelout<=1'b1;
15773: pixelout<=1'b1;
15774: pixelout<=1'b1;
15775: pixelout<=1'b1;
15776: pixelout<=1'b1;
15777: pixelout<=1'b1;
15778: pixelout<=1'b1;
15779: pixelout<=1'b1;
15780: pixelout<=1'b1;
15781: pixelout<=1'b1;
15782: pixelout<=1'b1;
15783: pixelout<=1'b1;
15784: pixelout<=1'b1;
15785: pixelout<=1'b1;
15786: pixelout<=1'b1;
15787: pixelout<=1'b1;
15788: pixelout<=1'b1;
15789: pixelout<=1'b1;
15790: pixelout<=1'b1;
15791: pixelout<=1'b1;
15792: pixelout<=1'b1;
15793: pixelout<=1'b1;
15794: pixelout<=1'b1;
15795: pixelout<=1'b1;
15796: pixelout<=1'b1;
15797: pixelout<=1'b1;
15798: pixelout<=1'b1;
15799: pixelout<=1'b1;
15800: pixelout<=1'b1;
15801: pixelout<=1'b1;
15802: pixelout<=1'b1;
15803: pixelout<=1'b1;
15804: pixelout<=1'b1;
15805: pixelout<=1'b1;
15806: pixelout<=1'b1;
15807: pixelout<=1'b1;
15808: pixelout<=1'b1;
15809: pixelout<=1'b1;
15810: pixelout<=1'b1;
15811: pixelout<=1'b1;
15812: pixelout<=1'b1;
15813: pixelout<=1'b1;
15814: pixelout<=1'b1;
15815: pixelout<=1'b1;
15816: pixelout<=1'b1;
15817: pixelout<=1'b1;
15818: pixelout<=1'b1;
15819: pixelout<=1'b1;
15820: pixelout<=1'b1;
15821: pixelout<=1'b1;
15822: pixelout<=1'b1;
15823: pixelout<=1'b1;
15824: pixelout<=1'b1;
15825: pixelout<=1'b1;
15826: pixelout<=1'b1;
15827: pixelout<=1'b1;
15828: pixelout<=1'b1;
15829: pixelout<=1'b1;
15830: pixelout<=1'b1;
15831: pixelout<=1'b1;
15832: pixelout<=1'b1;
15833: pixelout<=1'b1;
15834: pixelout<=1'b1;
15835: pixelout<=1'b1;
15836: pixelout<=1'b1;
15837: pixelout<=1'b1;
15838: pixelout<=1'b1;
15839: pixelout<=1'b1;
15840: pixelout<=1'b1;
15841: pixelout<=1'b1;
15842: pixelout<=1'b1;
15843: pixelout<=1'b1;
15844: pixelout<=1'b1;
15845: pixelout<=1'b1;
15846: pixelout<=1'b1;
15847: pixelout<=1'b1;
15848: pixelout<=1'b1;
15849: pixelout<=1'b1;
15850: pixelout<=1'b1;
15851: pixelout<=1'b1;
15852: pixelout<=1'b1;
15853: pixelout<=1'b1;
15854: pixelout<=1'b1;
15855: pixelout<=1'b1;
15856: pixelout<=1'b1;
15857: pixelout<=1'b1;
15858: pixelout<=1'b1;
15859: pixelout<=1'b1;
15860: pixelout<=1'b1;
15861: pixelout<=1'b1;
15862: pixelout<=1'b1;
15863: pixelout<=1'b1;
15864: pixelout<=1'b1;
15865: pixelout<=1'b1;
15866: pixelout<=1'b1;
15867: pixelout<=1'b1;
15868: pixelout<=1'b1;
15869: pixelout<=1'b1;
15870: pixelout<=1'b1;
15871: pixelout<=1'b1;
15872: pixelout<=1'b1;
15873: pixelout<=1'b1;
15874: pixelout<=1'b1;
15875: pixelout<=1'b1;
15876: pixelout<=1'b1;
15877: pixelout<=1'b1;
15878: pixelout<=1'b1;
15879: pixelout<=1'b1;
15880: pixelout<=1'b1;
15881: pixelout<=1'b1;
15882: pixelout<=1'b1;
15883: pixelout<=1'b1;
15884: pixelout<=1'b1;
15885: pixelout<=1'b1;
15886: pixelout<=1'b1;
15887: pixelout<=1'b1;
15888: pixelout<=1'b1;
15889: pixelout<=1'b1;
15890: pixelout<=1'b1;
15891: pixelout<=1'b1;
15892: pixelout<=1'b1;
15893: pixelout<=1'b1;
15894: pixelout<=1'b1;
15895: pixelout<=1'b1;
15896: pixelout<=1'b1;
15897: pixelout<=1'b1;
15898: pixelout<=1'b1;
15899: pixelout<=1'b1;
15900: pixelout<=1'b1;
15901: pixelout<=1'b1;
15902: pixelout<=1'b1;
15903: pixelout<=1'b1;
15904: pixelout<=1'b1;
15905: pixelout<=1'b1;
15906: pixelout<=1'b1;
15907: pixelout<=1'b1;
15908: pixelout<=1'b1;
15909: pixelout<=1'b1;
15910: pixelout<=1'b1;
15911: pixelout<=1'b1;
15912: pixelout<=1'b1;
15913: pixelout<=1'b1;
15914: pixelout<=1'b1;
15915: pixelout<=1'b1;
15916: pixelout<=1'b1;
15917: pixelout<=1'b1;
15918: pixelout<=1'b1;
15919: pixelout<=1'b1;
15920: pixelout<=1'b1;
15921: pixelout<=1'b1;
15922: pixelout<=1'b1;
15923: pixelout<=1'b1;
15924: pixelout<=1'b1;
15925: pixelout<=1'b1;
15926: pixelout<=1'b1;
15927: pixelout<=1'b1;
15928: pixelout<=1'b1;
15929: pixelout<=1'b1;
15930: pixelout<=1'b1;
15931: pixelout<=1'b1;
15932: pixelout<=1'b1;
15933: pixelout<=1'b1;
15934: pixelout<=1'b1;
15935: pixelout<=1'b1;
15936: pixelout<=1'b1;
15937: pixelout<=1'b1;
15938: pixelout<=1'b1;
15939: pixelout<=1'b1;
15940: pixelout<=1'b1;
15941: pixelout<=1'b1;
15942: pixelout<=1'b1;
15943: pixelout<=1'b1;
15944: pixelout<=1'b1;
15945: pixelout<=1'b1;
15946: pixelout<=1'b1;
15947: pixelout<=1'b1;
15948: pixelout<=1'b1;
15949: pixelout<=1'b1;
15950: pixelout<=1'b1;
15951: pixelout<=1'b1;
15952: pixelout<=1'b1;
15953: pixelout<=1'b1;
15954: pixelout<=1'b1;
15955: pixelout<=1'b1;
15956: pixelout<=1'b1;
15957: pixelout<=1'b1;
15958: pixelout<=1'b1;
15959: pixelout<=1'b1;
15960: pixelout<=1'b1;
15961: pixelout<=1'b1;
15962: pixelout<=1'b1;
15963: pixelout<=1'b1;
15964: pixelout<=1'b1;
15965: pixelout<=1'b1;
15966: pixelout<=1'b1;
15967: pixelout<=1'b1;
15968: pixelout<=1'b1;
15969: pixelout<=1'b1;
15970: pixelout<=1'b1;
15971: pixelout<=1'b1;
15972: pixelout<=1'b1;
15973: pixelout<=1'b1;
15974: pixelout<=1'b1;
15975: pixelout<=1'b1;
15976: pixelout<=1'b1;
15977: pixelout<=1'b1;
15978: pixelout<=1'b1;
15979: pixelout<=1'b1;
15980: pixelout<=1'b1;
15981: pixelout<=1'b1;
15982: pixelout<=1'b1;
15983: pixelout<=1'b1;
15984: pixelout<=1'b1;
15985: pixelout<=1'b1;
15986: pixelout<=1'b1;
15987: pixelout<=1'b1;
15988: pixelout<=1'b1;
15989: pixelout<=1'b1;
15990: pixelout<=1'b1;
15991: pixelout<=1'b1;
15992: pixelout<=1'b1;
15993: pixelout<=1'b1;
15994: pixelout<=1'b1;
15995: pixelout<=1'b1;
15996: pixelout<=1'b1;
15997: pixelout<=1'b1;
15998: pixelout<=1'b1;
15999: pixelout<=1'b1;
16000: pixelout<=1'b1;
16001: pixelout<=1'b1;
16002: pixelout<=1'b1;
16003: pixelout<=1'b1;
16004: pixelout<=1'b1;
16005: pixelout<=1'b1;
16006: pixelout<=1'b1;
16007: pixelout<=1'b1;
16008: pixelout<=1'b1;
16009: pixelout<=1'b1;
16010: pixelout<=1'b1;
16011: pixelout<=1'b1;
16012: pixelout<=1'b1;
16013: pixelout<=1'b1;
16014: pixelout<=1'b1;
16015: pixelout<=1'b1;
16016: pixelout<=1'b1;
16017: pixelout<=1'b1;
16018: pixelout<=1'b1;
16019: pixelout<=1'b1;
16020: pixelout<=1'b1;
16021: pixelout<=1'b1;
16022: pixelout<=1'b1;
16023: pixelout<=1'b1;
16024: pixelout<=1'b1;
16025: pixelout<=1'b1;
16026: pixelout<=1'b1;
16027: pixelout<=1'b1;
16028: pixelout<=1'b1;
16029: pixelout<=1'b1;
16030: pixelout<=1'b1;
16031: pixelout<=1'b1;
16032: pixelout<=1'b1;
16033: pixelout<=1'b1;
16034: pixelout<=1'b1;
16035: pixelout<=1'b1;
16036: pixelout<=1'b1;
16037: pixelout<=1'b1;
16038: pixelout<=1'b1;
16039: pixelout<=1'b1;
16040: pixelout<=1'b1;
16041: pixelout<=1'b1;
16042: pixelout<=1'b1;
16043: pixelout<=1'b1;
16044: pixelout<=1'b1;
16045: pixelout<=1'b1;
16046: pixelout<=1'b1;
16047: pixelout<=1'b1;
16048: pixelout<=1'b1;
16049: pixelout<=1'b1;
16050: pixelout<=1'b1;
16051: pixelout<=1'b1;
16052: pixelout<=1'b1;
16053: pixelout<=1'b1;
16054: pixelout<=1'b1;
16055: pixelout<=1'b1;
16056: pixelout<=1'b1;
16057: pixelout<=1'b1;
16058: pixelout<=1'b1;
16059: pixelout<=1'b1;
16060: pixelout<=1'b1;
16061: pixelout<=1'b1;
16062: pixelout<=1'b1;
16063: pixelout<=1'b1;
16064: pixelout<=1'b1;
16065: pixelout<=1'b1;
16066: pixelout<=1'b1;
16067: pixelout<=1'b1;
16068: pixelout<=1'b1;
16069: pixelout<=1'b1;
16070: pixelout<=1'b1;
16071: pixelout<=1'b1;
16072: pixelout<=1'b1;
16073: pixelout<=1'b1;
16074: pixelout<=1'b1;
16075: pixelout<=1'b1;
16076: pixelout<=1'b1;
16077: pixelout<=1'b1;
16078: pixelout<=1'b1;
16079: pixelout<=1'b1;
16080: pixelout<=1'b1;
16081: pixelout<=1'b1;
16082: pixelout<=1'b1;
16083: pixelout<=1'b1;
16084: pixelout<=1'b1;
16085: pixelout<=1'b1;
16086: pixelout<=1'b1;
16087: pixelout<=1'b1;
16088: pixelout<=1'b1;
16089: pixelout<=1'b1;
16090: pixelout<=1'b1;
16091: pixelout<=1'b1;
16092: pixelout<=1'b1;
16093: pixelout<=1'b1;
16094: pixelout<=1'b1;
16095: pixelout<=1'b1;
16096: pixelout<=1'b1;
16097: pixelout<=1'b1;
16098: pixelout<=1'b1;
16099: pixelout<=1'b1;
16100: pixelout<=1'b1;
16101: pixelout<=1'b1;
16102: pixelout<=1'b1;
16103: pixelout<=1'b1;
16104: pixelout<=1'b1;
16105: pixelout<=1'b1;
16106: pixelout<=1'b1;
16107: pixelout<=1'b1;
16108: pixelout<=1'b1;
16109: pixelout<=1'b1;
16110: pixelout<=1'b1;
16111: pixelout<=1'b1;
16112: pixelout<=1'b1;
16113: pixelout<=1'b1;
16114: pixelout<=1'b1;
16115: pixelout<=1'b1;
16116: pixelout<=1'b1;
16117: pixelout<=1'b1;
16118: pixelout<=1'b1;
16119: pixelout<=1'b1;
16120: pixelout<=1'b1;
16121: pixelout<=1'b1;
16122: pixelout<=1'b1;
16123: pixelout<=1'b1;
16124: pixelout<=1'b1;
16125: pixelout<=1'b1;
16126: pixelout<=1'b1;
16127: pixelout<=1'b1;
16128: pixelout<=1'b1;
16129: pixelout<=1'b1;
16130: pixelout<=1'b1;
16131: pixelout<=1'b1;
16132: pixelout<=1'b1;
16133: pixelout<=1'b1;
16134: pixelout<=1'b1;
16135: pixelout<=1'b1;
16136: pixelout<=1'b1;
16137: pixelout<=1'b1;
16138: pixelout<=1'b1;
16139: pixelout<=1'b1;
16140: pixelout<=1'b1;
16141: pixelout<=1'b1;
16142: pixelout<=1'b1;
16143: pixelout<=1'b1;
16144: pixelout<=1'b1;
16145: pixelout<=1'b1;
16146: pixelout<=1'b1;
16147: pixelout<=1'b1;
16148: pixelout<=1'b1;
16149: pixelout<=1'b1;
16150: pixelout<=1'b1;
16151: pixelout<=1'b1;
16152: pixelout<=1'b1;
16153: pixelout<=1'b1;
16154: pixelout<=1'b1;
16155: pixelout<=1'b1;
16156: pixelout<=1'b1;
16157: pixelout<=1'b1;
16158: pixelout<=1'b1;
16159: pixelout<=1'b1;
16160: pixelout<=1'b1;
16161: pixelout<=1'b1;
16162: pixelout<=1'b1;
16163: pixelout<=1'b1;
16164: pixelout<=1'b1;
16165: pixelout<=1'b1;
16166: pixelout<=1'b1;
16167: pixelout<=1'b1;
16168: pixelout<=1'b1;
16169: pixelout<=1'b1;
16170: pixelout<=1'b1;
16171: pixelout<=1'b1;
16172: pixelout<=1'b1;
16173: pixelout<=1'b1;
16174: pixelout<=1'b1;
16175: pixelout<=1'b1;
16176: pixelout<=1'b1;
16177: pixelout<=1'b1;
16178: pixelout<=1'b1;
16179: pixelout<=1'b1;
16180: pixelout<=1'b1;
16181: pixelout<=1'b1;
16182: pixelout<=1'b1;
16183: pixelout<=1'b1;
16184: pixelout<=1'b1;
16185: pixelout<=1'b1;
16186: pixelout<=1'b1;
16187: pixelout<=1'b1;
16188: pixelout<=1'b1;
16189: pixelout<=1'b1;
16190: pixelout<=1'b1;
16191: pixelout<=1'b1;
16192: pixelout<=1'b1;
16193: pixelout<=1'b1;
16194: pixelout<=1'b1;
16195: pixelout<=1'b1;
16196: pixelout<=1'b1;
16197: pixelout<=1'b1;
16198: pixelout<=1'b1;
16199: pixelout<=1'b1;
16200: pixelout<=1'b1;
16201: pixelout<=1'b1;
16202: pixelout<=1'b1;
16203: pixelout<=1'b1;
16204: pixelout<=1'b1;
16205: pixelout<=1'b1;
16206: pixelout<=1'b1;
16207: pixelout<=1'b1;
16208: pixelout<=1'b1;
16209: pixelout<=1'b1;
16210: pixelout<=1'b1;
16211: pixelout<=1'b1;
16212: pixelout<=1'b1;
16213: pixelout<=1'b1;
16214: pixelout<=1'b1;
16215: pixelout<=1'b1;
16216: pixelout<=1'b1;
16217: pixelout<=1'b1;
16218: pixelout<=1'b1;
16219: pixelout<=1'b1;
16220: pixelout<=1'b1;
16221: pixelout<=1'b1;
16222: pixelout<=1'b1;
16223: pixelout<=1'b1;
16224: pixelout<=1'b1;
16225: pixelout<=1'b1;
16226: pixelout<=1'b1;
16227: pixelout<=1'b1;
16228: pixelout<=1'b1;
16229: pixelout<=1'b1;
16230: pixelout<=1'b1;
16231: pixelout<=1'b1;
16232: pixelout<=1'b1;
16233: pixelout<=1'b1;
16234: pixelout<=1'b1;
16235: pixelout<=1'b1;
16236: pixelout<=1'b1;
16237: pixelout<=1'b1;
16238: pixelout<=1'b1;
16239: pixelout<=1'b1;
16240: pixelout<=1'b1;
16241: pixelout<=1'b1;
16242: pixelout<=1'b1;
16243: pixelout<=1'b1;
16244: pixelout<=1'b1;
16245: pixelout<=1'b1;
16246: pixelout<=1'b1;
16247: pixelout<=1'b1;
16248: pixelout<=1'b1;
16249: pixelout<=1'b1;
16250: pixelout<=1'b1;
16251: pixelout<=1'b1;
16252: pixelout<=1'b1;
16253: pixelout<=1'b1;
16254: pixelout<=1'b1;
16255: pixelout<=1'b1;
16256: pixelout<=1'b1;
16257: pixelout<=1'b1;
16258: pixelout<=1'b1;
16259: pixelout<=1'b1;
16260: pixelout<=1'b1;
16261: pixelout<=1'b1;
16262: pixelout<=1'b1;
16263: pixelout<=1'b1;
16264: pixelout<=1'b1;
16265: pixelout<=1'b1;
16266: pixelout<=1'b1;
16267: pixelout<=1'b1;
16268: pixelout<=1'b1;
16269: pixelout<=1'b1;
16270: pixelout<=1'b1;
16271: pixelout<=1'b1;
16272: pixelout<=1'b1;
16273: pixelout<=1'b1;
16274: pixelout<=1'b1;
16275: pixelout<=1'b1;
16276: pixelout<=1'b1;
16277: pixelout<=1'b1;
16278: pixelout<=1'b1;
16279: pixelout<=1'b1;
16280: pixelout<=1'b1;
16281: pixelout<=1'b1;
16282: pixelout<=1'b1;
16283: pixelout<=1'b1;
16284: pixelout<=1'b1;
16285: pixelout<=1'b1;
16286: pixelout<=1'b1;
16287: pixelout<=1'b1;
16288: pixelout<=1'b1;
16289: pixelout<=1'b1;
16290: pixelout<=1'b1;
16291: pixelout<=1'b1;
16292: pixelout<=1'b1;
16293: pixelout<=1'b1;
16294: pixelout<=1'b1;
16295: pixelout<=1'b1;
16296: pixelout<=1'b1;
16297: pixelout<=1'b1;
16298: pixelout<=1'b1;
16299: pixelout<=1'b1;
16300: pixelout<=1'b1;
16301: pixelout<=1'b1;
16302: pixelout<=1'b1;
16303: pixelout<=1'b1;
16304: pixelout<=1'b1;
16305: pixelout<=1'b1;
16306: pixelout<=1'b1;
16307: pixelout<=1'b1;
16308: pixelout<=1'b1;
16309: pixelout<=1'b1;
16310: pixelout<=1'b1;
16311: pixelout<=1'b1;
16312: pixelout<=1'b1;
16313: pixelout<=1'b1;
16314: pixelout<=1'b1;
16315: pixelout<=1'b1;
16316: pixelout<=1'b1;
16317: pixelout<=1'b1;
16318: pixelout<=1'b1;
16319: pixelout<=1'b1;
16320: pixelout<=1'b1;
16321: pixelout<=1'b1;
16322: pixelout<=1'b1;
16323: pixelout<=1'b1;
16324: pixelout<=1'b1;
16325: pixelout<=1'b1;
16326: pixelout<=1'b1;
16327: pixelout<=1'b1;
16328: pixelout<=1'b1;
16329: pixelout<=1'b1;
16330: pixelout<=1'b1;
16331: pixelout<=1'b1;
16332: pixelout<=1'b1;
16333: pixelout<=1'b1;
16334: pixelout<=1'b1;
16335: pixelout<=1'b1;
16336: pixelout<=1'b1;
16337: pixelout<=1'b1;
16338: pixelout<=1'b1;
16339: pixelout<=1'b1;
16340: pixelout<=1'b1;
16341: pixelout<=1'b1;
16342: pixelout<=1'b1;
16343: pixelout<=1'b1;
16344: pixelout<=1'b1;
16345: pixelout<=1'b1;
16346: pixelout<=1'b1;
16347: pixelout<=1'b1;
16348: pixelout<=1'b1;
16349: pixelout<=1'b1;
16350: pixelout<=1'b1;
16351: pixelout<=1'b1;
16352: pixelout<=1'b1;
16353: pixelout<=1'b1;
16354: pixelout<=1'b1;
16355: pixelout<=1'b1;
16356: pixelout<=1'b1;
16357: pixelout<=1'b1;
16358: pixelout<=1'b1;
16359: pixelout<=1'b1;
16360: pixelout<=1'b1;
16361: pixelout<=1'b1;
16362: pixelout<=1'b1;
16363: pixelout<=1'b1;
16364: pixelout<=1'b1;
16365: pixelout<=1'b1;
16366: pixelout<=1'b1;
16367: pixelout<=1'b1;
16368: pixelout<=1'b1;
16369: pixelout<=1'b1;
16370: pixelout<=1'b1;
16371: pixelout<=1'b1;
16372: pixelout<=1'b1;
16373: pixelout<=1'b1;
16374: pixelout<=1'b1;
16375: pixelout<=1'b1;
16376: pixelout<=1'b1;
16377: pixelout<=1'b1;
16378: pixelout<=1'b1;
16379: pixelout<=1'b1;
16380: pixelout<=1'b1;
16381: pixelout<=1'b1;
16382: pixelout<=1'b1;
16383: pixelout<=1'b1;
16384: pixelout<=1'b1;
16385: pixelout<=1'b1;
16386: pixelout<=1'b1;
16387: pixelout<=1'b1;
16388: pixelout<=1'b1;
16389: pixelout<=1'b1;
16390: pixelout<=1'b1;
16391: pixelout<=1'b1;
16392: pixelout<=1'b1;
16393: pixelout<=1'b1;
16394: pixelout<=1'b1;
16395: pixelout<=1'b1;
16396: pixelout<=1'b1;
16397: pixelout<=1'b1;
16398: pixelout<=1'b1;
16399: pixelout<=1'b1;
16400: pixelout<=1'b1;
16401: pixelout<=1'b1;
16402: pixelout<=1'b1;
16403: pixelout<=1'b1;
16404: pixelout<=1'b1;
16405: pixelout<=1'b1;
16406: pixelout<=1'b1;
16407: pixelout<=1'b1;
16408: pixelout<=1'b1;
16409: pixelout<=1'b1;
16410: pixelout<=1'b1;
16411: pixelout<=1'b1;
16412: pixelout<=1'b1;
16413: pixelout<=1'b1;
16414: pixelout<=1'b1;
16415: pixelout<=1'b1;
16416: pixelout<=1'b1;
16417: pixelout<=1'b1;
16418: pixelout<=1'b1;
16419: pixelout<=1'b1;
16420: pixelout<=1'b1;
16421: pixelout<=1'b1;
16422: pixelout<=1'b1;
16423: pixelout<=1'b1;
16424: pixelout<=1'b1;
16425: pixelout<=1'b1;
16426: pixelout<=1'b1;
16427: pixelout<=1'b1;
16428: pixelout<=1'b1;
16429: pixelout<=1'b1;
16430: pixelout<=1'b1;
16431: pixelout<=1'b1;
16432: pixelout<=1'b1;
16433: pixelout<=1'b1;
16434: pixelout<=1'b1;
16435: pixelout<=1'b1;
16436: pixelout<=1'b1;
16437: pixelout<=1'b1;
16438: pixelout<=1'b1;
16439: pixelout<=1'b1;
16440: pixelout<=1'b1;
16441: pixelout<=1'b1;
16442: pixelout<=1'b1;
16443: pixelout<=1'b1;
16444: pixelout<=1'b1;
16445: pixelout<=1'b1;
16446: pixelout<=1'b1;
16447: pixelout<=1'b1;
16448: pixelout<=1'b1;
16449: pixelout<=1'b1;
16450: pixelout<=1'b1;
16451: pixelout<=1'b1;
16452: pixelout<=1'b1;
16453: pixelout<=1'b1;
16454: pixelout<=1'b1;
16455: pixelout<=1'b1;
16456: pixelout<=1'b1;
16457: pixelout<=1'b1;
16458: pixelout<=1'b1;
16459: pixelout<=1'b1;
16460: pixelout<=1'b1;
16461: pixelout<=1'b1;
16462: pixelout<=1'b1;
16463: pixelout<=1'b1;
16464: pixelout<=1'b1;
16465: pixelout<=1'b1;
16466: pixelout<=1'b1;
16467: pixelout<=1'b1;
16468: pixelout<=1'b1;
16469: pixelout<=1'b1;
16470: pixelout<=1'b1;
16471: pixelout<=1'b1;
16472: pixelout<=1'b1;
16473: pixelout<=1'b1;
16474: pixelout<=1'b1;
16475: pixelout<=1'b1;
16476: pixelout<=1'b1;
16477: pixelout<=1'b1;
16478: pixelout<=1'b1;
16479: pixelout<=1'b1;
16480: pixelout<=1'b1;
16481: pixelout<=1'b1;
16482: pixelout<=1'b1;
16483: pixelout<=1'b1;
16484: pixelout<=1'b1;
16485: pixelout<=1'b1;
16486: pixelout<=1'b1;
16487: pixelout<=1'b1;
16488: pixelout<=1'b1;
16489: pixelout<=1'b1;
16490: pixelout<=1'b1;
16491: pixelout<=1'b1;
16492: pixelout<=1'b1;
16493: pixelout<=1'b1;
16494: pixelout<=1'b1;
16495: pixelout<=1'b1;
16496: pixelout<=1'b1;
16497: pixelout<=1'b1;
16498: pixelout<=1'b1;
16499: pixelout<=1'b1;
16500: pixelout<=1'b1;
16501: pixelout<=1'b1;
16502: pixelout<=1'b1;
16503: pixelout<=1'b1;
16504: pixelout<=1'b1;
16505: pixelout<=1'b1;
16506: pixelout<=1'b1;
16507: pixelout<=1'b1;
16508: pixelout<=1'b1;
16509: pixelout<=1'b1;
16510: pixelout<=1'b1;
16511: pixelout<=1'b1;
16512: pixelout<=1'b1;
16513: pixelout<=1'b1;
16514: pixelout<=1'b1;
16515: pixelout<=1'b1;
16516: pixelout<=1'b1;
16517: pixelout<=1'b1;
16518: pixelout<=1'b1;
16519: pixelout<=1'b1;
16520: pixelout<=1'b1;
16521: pixelout<=1'b1;
16522: pixelout<=1'b1;
16523: pixelout<=1'b1;
16524: pixelout<=1'b1;
16525: pixelout<=1'b1;
16526: pixelout<=1'b1;
16527: pixelout<=1'b1;
16528: pixelout<=1'b1;
16529: pixelout<=1'b1;
16530: pixelout<=1'b1;
16531: pixelout<=1'b1;
16532: pixelout<=1'b1;
16533: pixelout<=1'b1;
16534: pixelout<=1'b1;
16535: pixelout<=1'b1;
16536: pixelout<=1'b1;
16537: pixelout<=1'b1;
16538: pixelout<=1'b1;
16539: pixelout<=1'b1;
16540: pixelout<=1'b1;
16541: pixelout<=1'b1;
16542: pixelout<=1'b1;
16543: pixelout<=1'b1;
16544: pixelout<=1'b1;
16545: pixelout<=1'b1;
16546: pixelout<=1'b1;
16547: pixelout<=1'b1;
16548: pixelout<=1'b1;
16549: pixelout<=1'b1;
16550: pixelout<=1'b1;
16551: pixelout<=1'b1;
16552: pixelout<=1'b1;
16553: pixelout<=1'b1;
16554: pixelout<=1'b1;
16555: pixelout<=1'b1;
16556: pixelout<=1'b1;
16557: pixelout<=1'b1;
16558: pixelout<=1'b1;
16559: pixelout<=1'b1;
16560: pixelout<=1'b1;
16561: pixelout<=1'b1;
16562: pixelout<=1'b1;
16563: pixelout<=1'b1;
16564: pixelout<=1'b1;
16565: pixelout<=1'b1;
16566: pixelout<=1'b1;
16567: pixelout<=1'b1;
16568: pixelout<=1'b1;
16569: pixelout<=1'b1;
16570: pixelout<=1'b1;
16571: pixelout<=1'b1;
16572: pixelout<=1'b1;
16573: pixelout<=1'b1;
16574: pixelout<=1'b1;
16575: pixelout<=1'b1;
16576: pixelout<=1'b1;
16577: pixelout<=1'b1;
16578: pixelout<=1'b1;
16579: pixelout<=1'b1;
16580: pixelout<=1'b1;
16581: pixelout<=1'b1;
16582: pixelout<=1'b1;
16583: pixelout<=1'b1;
16584: pixelout<=1'b1;
16585: pixelout<=1'b1;
16586: pixelout<=1'b1;
16587: pixelout<=1'b1;
16588: pixelout<=1'b1;
16589: pixelout<=1'b1;
16590: pixelout<=1'b1;
16591: pixelout<=1'b1;
16592: pixelout<=1'b1;
16593: pixelout<=1'b1;
16594: pixelout<=1'b1;
16595: pixelout<=1'b1;
16596: pixelout<=1'b1;
16597: pixelout<=1'b1;
16598: pixelout<=1'b1;
16599: pixelout<=1'b1;
16600: pixelout<=1'b1;
16601: pixelout<=1'b1;
16602: pixelout<=1'b1;
16603: pixelout<=1'b1;
16604: pixelout<=1'b1;
16605: pixelout<=1'b1;
16606: pixelout<=1'b1;
16607: pixelout<=1'b1;
16608: pixelout<=1'b1;
16609: pixelout<=1'b1;
16610: pixelout<=1'b1;
16611: pixelout<=1'b1;
16612: pixelout<=1'b1;
16613: pixelout<=1'b1;
16614: pixelout<=1'b1;
16615: pixelout<=1'b1;
16616: pixelout<=1'b1;
16617: pixelout<=1'b1;
16618: pixelout<=1'b1;
16619: pixelout<=1'b1;
16620: pixelout<=1'b1;
16621: pixelout<=1'b1;
16622: pixelout<=1'b1;
16623: pixelout<=1'b1;
16624: pixelout<=1'b1;
16625: pixelout<=1'b1;
16626: pixelout<=1'b1;
16627: pixelout<=1'b1;
16628: pixelout<=1'b1;
16629: pixelout<=1'b1;
16630: pixelout<=1'b1;
16631: pixelout<=1'b1;
16632: pixelout<=1'b1;
16633: pixelout<=1'b1;
16634: pixelout<=1'b1;
16635: pixelout<=1'b1;
16636: pixelout<=1'b1;
16637: pixelout<=1'b1;
16638: pixelout<=1'b1;
16639: pixelout<=1'b1;
16640: pixelout<=1'b1;
16641: pixelout<=1'b1;
16642: pixelout<=1'b1;
16643: pixelout<=1'b1;
16644: pixelout<=1'b1;
16645: pixelout<=1'b1;
16646: pixelout<=1'b1;
16647: pixelout<=1'b1;
16648: pixelout<=1'b1;
16649: pixelout<=1'b1;
16650: pixelout<=1'b1;
16651: pixelout<=1'b1;
16652: pixelout<=1'b1;
16653: pixelout<=1'b1;
16654: pixelout<=1'b1;
16655: pixelout<=1'b1;
16656: pixelout<=1'b1;
16657: pixelout<=1'b1;
16658: pixelout<=1'b1;
16659: pixelout<=1'b1;
16660: pixelout<=1'b1;
16661: pixelout<=1'b1;
16662: pixelout<=1'b1;
16663: pixelout<=1'b1;
16664: pixelout<=1'b1;
16665: pixelout<=1'b1;
16666: pixelout<=1'b1;
16667: pixelout<=1'b1;
16668: pixelout<=1'b1;
16669: pixelout<=1'b1;
16670: pixelout<=1'b1;
16671: pixelout<=1'b1;
16672: pixelout<=1'b1;
16673: pixelout<=1'b1;
16674: pixelout<=1'b1;
16675: pixelout<=1'b1;
16676: pixelout<=1'b1;
16677: pixelout<=1'b1;
16678: pixelout<=1'b1;
16679: pixelout<=1'b1;
16680: pixelout<=1'b1;
16681: pixelout<=1'b1;
16682: pixelout<=1'b1;
16683: pixelout<=1'b1;
16684: pixelout<=1'b1;
16685: pixelout<=1'b1;
16686: pixelout<=1'b1;
16687: pixelout<=1'b1;
16688: pixelout<=1'b1;
16689: pixelout<=1'b1;
16690: pixelout<=1'b1;
16691: pixelout<=1'b1;
16692: pixelout<=1'b1;
16693: pixelout<=1'b1;
16694: pixelout<=1'b1;
16695: pixelout<=1'b1;
16696: pixelout<=1'b1;
16697: pixelout<=1'b1;
16698: pixelout<=1'b1;
16699: pixelout<=1'b1;
16700: pixelout<=1'b1;
16701: pixelout<=1'b1;
16702: pixelout<=1'b1;
16703: pixelout<=1'b1;
16704: pixelout<=1'b1;
16705: pixelout<=1'b1;
16706: pixelout<=1'b1;
16707: pixelout<=1'b1;
16708: pixelout<=1'b1;
16709: pixelout<=1'b1;
16710: pixelout<=1'b1;
16711: pixelout<=1'b1;
16712: pixelout<=1'b1;
16713: pixelout<=1'b1;
16714: pixelout<=1'b1;
16715: pixelout<=1'b1;
16716: pixelout<=1'b1;
16717: pixelout<=1'b1;
16718: pixelout<=1'b1;
16719: pixelout<=1'b1;
16720: pixelout<=1'b1;
16721: pixelout<=1'b1;
16722: pixelout<=1'b1;
16723: pixelout<=1'b1;
16724: pixelout<=1'b1;
16725: pixelout<=1'b1;
16726: pixelout<=1'b1;
16727: pixelout<=1'b1;
16728: pixelout<=1'b1;
16729: pixelout<=1'b1;
16730: pixelout<=1'b1;
16731: pixelout<=1'b1;
16732: pixelout<=1'b1;
16733: pixelout<=1'b1;
16734: pixelout<=1'b1;
16735: pixelout<=1'b1;
16736: pixelout<=1'b1;
16737: pixelout<=1'b1;
16738: pixelout<=1'b1;
16739: pixelout<=1'b1;
16740: pixelout<=1'b1;
16741: pixelout<=1'b1;
16742: pixelout<=1'b1;
16743: pixelout<=1'b1;
16744: pixelout<=1'b1;
16745: pixelout<=1'b1;
16746: pixelout<=1'b1;
16747: pixelout<=1'b1;
16748: pixelout<=1'b1;
16749: pixelout<=1'b1;
16750: pixelout<=1'b1;
16751: pixelout<=1'b1;
16752: pixelout<=1'b1;
16753: pixelout<=1'b1;
16754: pixelout<=1'b1;
16755: pixelout<=1'b1;
16756: pixelout<=1'b1;
16757: pixelout<=1'b1;
16758: pixelout<=1'b1;
16759: pixelout<=1'b1;
16760: pixelout<=1'b1;
16761: pixelout<=1'b1;
16762: pixelout<=1'b1;
16763: pixelout<=1'b1;
16764: pixelout<=1'b1;
16765: pixelout<=1'b1;
16766: pixelout<=1'b1;
16767: pixelout<=1'b1;
16768: pixelout<=1'b1;
16769: pixelout<=1'b1;
16770: pixelout<=1'b1;
16771: pixelout<=1'b1;
16772: pixelout<=1'b1;
16773: pixelout<=1'b1;
16774: pixelout<=1'b1;
16775: pixelout<=1'b1;
16776: pixelout<=1'b1;
16777: pixelout<=1'b1;
16778: pixelout<=1'b1;
16779: pixelout<=1'b1;
16780: pixelout<=1'b1;
16781: pixelout<=1'b1;
16782: pixelout<=1'b1;
16783: pixelout<=1'b1;
16784: pixelout<=1'b1;
16785: pixelout<=1'b1;
16786: pixelout<=1'b1;
16787: pixelout<=1'b1;
16788: pixelout<=1'b1;
16789: pixelout<=1'b1;
16790: pixelout<=1'b1;
16791: pixelout<=1'b1;
16792: pixelout<=1'b1;
16793: pixelout<=1'b1;
16794: pixelout<=1'b1;
16795: pixelout<=1'b1;
16796: pixelout<=1'b1;
16797: pixelout<=1'b1;
16798: pixelout<=1'b1;
16799: pixelout<=1'b1;
16800: pixelout<=1'b1;
16801: pixelout<=1'b1;
16802: pixelout<=1'b1;
16803: pixelout<=1'b1;
16804: pixelout<=1'b1;
16805: pixelout<=1'b1;
16806: pixelout<=1'b1;
16807: pixelout<=1'b1;
16808: pixelout<=1'b1;
16809: pixelout<=1'b1;
16810: pixelout<=1'b1;
16811: pixelout<=1'b1;
16812: pixelout<=1'b1;
16813: pixelout<=1'b1;
16814: pixelout<=1'b1;
16815: pixelout<=1'b1;
16816: pixelout<=1'b1;
16817: pixelout<=1'b1;
16818: pixelout<=1'b1;
16819: pixelout<=1'b1;
16820: pixelout<=1'b1;
16821: pixelout<=1'b1;
16822: pixelout<=1'b1;
16823: pixelout<=1'b1;
16824: pixelout<=1'b1;
16825: pixelout<=1'b1;
16826: pixelout<=1'b1;
16827: pixelout<=1'b1;
16828: pixelout<=1'b1;
16829: pixelout<=1'b1;
16830: pixelout<=1'b1;
16831: pixelout<=1'b1;
16832: pixelout<=1'b1;
16833: pixelout<=1'b1;
16834: pixelout<=1'b1;
16835: pixelout<=1'b1;
16836: pixelout<=1'b1;
16837: pixelout<=1'b1;
16838: pixelout<=1'b1;
16839: pixelout<=1'b1;
16840: pixelout<=1'b1;
16841: pixelout<=1'b1;
16842: pixelout<=1'b1;
16843: pixelout<=1'b1;
16844: pixelout<=1'b1;
16845: pixelout<=1'b1;
16846: pixelout<=1'b1;
16847: pixelout<=1'b1;
16848: pixelout<=1'b1;
16849: pixelout<=1'b1;
16850: pixelout<=1'b1;
16851: pixelout<=1'b1;
16852: pixelout<=1'b1;
16853: pixelout<=1'b1;
16854: pixelout<=1'b1;
16855: pixelout<=1'b1;
16856: pixelout<=1'b1;
16857: pixelout<=1'b1;
16858: pixelout<=1'b1;
16859: pixelout<=1'b1;
16860: pixelout<=1'b1;
16861: pixelout<=1'b1;
16862: pixelout<=1'b1;
16863: pixelout<=1'b1;
16864: pixelout<=1'b1;
16865: pixelout<=1'b1;
16866: pixelout<=1'b1;
16867: pixelout<=1'b1;
16868: pixelout<=1'b1;
16869: pixelout<=1'b1;
16870: pixelout<=1'b1;
16871: pixelout<=1'b1;
16872: pixelout<=1'b1;
16873: pixelout<=1'b1;
16874: pixelout<=1'b1;
16875: pixelout<=1'b1;
16876: pixelout<=1'b1;
16877: pixelout<=1'b1;
16878: pixelout<=1'b1;
16879: pixelout<=1'b1;
16880: pixelout<=1'b1;
16881: pixelout<=1'b1;
16882: pixelout<=1'b1;
16883: pixelout<=1'b1;
16884: pixelout<=1'b1;
16885: pixelout<=1'b1;
16886: pixelout<=1'b1;
16887: pixelout<=1'b1;
16888: pixelout<=1'b1;
16889: pixelout<=1'b1;
16890: pixelout<=1'b1;
16891: pixelout<=1'b1;
16892: pixelout<=1'b1;
16893: pixelout<=1'b1;
16894: pixelout<=1'b1;
16895: pixelout<=1'b1;
16896: pixelout<=1'b1;
16897: pixelout<=1'b1;
16898: pixelout<=1'b1;
16899: pixelout<=1'b1;
16900: pixelout<=1'b1;
16901: pixelout<=1'b1;
16902: pixelout<=1'b1;
16903: pixelout<=1'b1;
16904: pixelout<=1'b1;
16905: pixelout<=1'b1;
16906: pixelout<=1'b1;
16907: pixelout<=1'b1;
16908: pixelout<=1'b1;
16909: pixelout<=1'b1;
16910: pixelout<=1'b1;
16911: pixelout<=1'b1;
16912: pixelout<=1'b1;
16913: pixelout<=1'b1;
16914: pixelout<=1'b1;
16915: pixelout<=1'b1;
16916: pixelout<=1'b1;
16917: pixelout<=1'b1;
16918: pixelout<=1'b1;
16919: pixelout<=1'b1;
16920: pixelout<=1'b1;
16921: pixelout<=1'b1;
16922: pixelout<=1'b1;
16923: pixelout<=1'b1;
16924: pixelout<=1'b1;
16925: pixelout<=1'b1;
16926: pixelout<=1'b1;
16927: pixelout<=1'b1;
16928: pixelout<=1'b1;
16929: pixelout<=1'b1;
16930: pixelout<=1'b1;
16931: pixelout<=1'b1;
16932: pixelout<=1'b1;
16933: pixelout<=1'b1;
16934: pixelout<=1'b1;
16935: pixelout<=1'b1;
16936: pixelout<=1'b1;
16937: pixelout<=1'b1;
16938: pixelout<=1'b1;
16939: pixelout<=1'b1;
16940: pixelout<=1'b1;
16941: pixelout<=1'b1;
16942: pixelout<=1'b1;
16943: pixelout<=1'b1;
16944: pixelout<=1'b1;
16945: pixelout<=1'b1;
16946: pixelout<=1'b1;
16947: pixelout<=1'b1;
16948: pixelout<=1'b1;
16949: pixelout<=1'b1;
16950: pixelout<=1'b1;
16951: pixelout<=1'b1;
16952: pixelout<=1'b1;
16953: pixelout<=1'b1;
16954: pixelout<=1'b1;
16955: pixelout<=1'b1;
16956: pixelout<=1'b1;
16957: pixelout<=1'b1;
16958: pixelout<=1'b1;
16959: pixelout<=1'b1;
16960: pixelout<=1'b1;
16961: pixelout<=1'b1;
16962: pixelout<=1'b1;
16963: pixelout<=1'b1;
16964: pixelout<=1'b1;
16965: pixelout<=1'b1;
16966: pixelout<=1'b1;
16967: pixelout<=1'b1;
16968: pixelout<=1'b1;
16969: pixelout<=1'b1;
16970: pixelout<=1'b1;
16971: pixelout<=1'b1;
16972: pixelout<=1'b1;
16973: pixelout<=1'b1;
16974: pixelout<=1'b1;
16975: pixelout<=1'b1;
16976: pixelout<=1'b1;
16977: pixelout<=1'b1;
16978: pixelout<=1'b1;
16979: pixelout<=1'b1;
16980: pixelout<=1'b1;
16981: pixelout<=1'b1;
16982: pixelout<=1'b1;
16983: pixelout<=1'b1;
16984: pixelout<=1'b1;
16985: pixelout<=1'b1;
16986: pixelout<=1'b1;
16987: pixelout<=1'b1;
16988: pixelout<=1'b1;
16989: pixelout<=1'b1;
16990: pixelout<=1'b1;
16991: pixelout<=1'b1;
16992: pixelout<=1'b1;
16993: pixelout<=1'b1;
16994: pixelout<=1'b1;
16995: pixelout<=1'b1;
16996: pixelout<=1'b1;
16997: pixelout<=1'b1;
16998: pixelout<=1'b1;
16999: pixelout<=1'b1;
17000: pixelout<=1'b1;
17001: pixelout<=1'b1;
17002: pixelout<=1'b1;
17003: pixelout<=1'b1;
17004: pixelout<=1'b1;
17005: pixelout<=1'b1;
17006: pixelout<=1'b1;
17007: pixelout<=1'b1;
17008: pixelout<=1'b1;
17009: pixelout<=1'b1;
17010: pixelout<=1'b1;
17011: pixelout<=1'b1;
17012: pixelout<=1'b1;
17013: pixelout<=1'b1;
17014: pixelout<=1'b1;
17015: pixelout<=1'b1;
17016: pixelout<=1'b1;
17017: pixelout<=1'b1;
17018: pixelout<=1'b1;
17019: pixelout<=1'b1;
17020: pixelout<=1'b1;
17021: pixelout<=1'b1;
17022: pixelout<=1'b1;
17023: pixelout<=1'b1;
17024: pixelout<=1'b1;
17025: pixelout<=1'b1;
17026: pixelout<=1'b1;
17027: pixelout<=1'b1;
17028: pixelout<=1'b1;
17029: pixelout<=1'b1;
17030: pixelout<=1'b1;
17031: pixelout<=1'b1;
17032: pixelout<=1'b1;
17033: pixelout<=1'b1;
17034: pixelout<=1'b1;
17035: pixelout<=1'b1;
17036: pixelout<=1'b1;
17037: pixelout<=1'b1;
17038: pixelout<=1'b1;
17039: pixelout<=1'b1;
17040: pixelout<=1'b1;
17041: pixelout<=1'b1;
17042: pixelout<=1'b1;
17043: pixelout<=1'b1;
17044: pixelout<=1'b1;
17045: pixelout<=1'b1;
17046: pixelout<=1'b1;
17047: pixelout<=1'b1;
17048: pixelout<=1'b1;
17049: pixelout<=1'b1;
17050: pixelout<=1'b0;
17051: pixelout<=1'b0;
17052: pixelout<=1'b0;
17053: pixelout<=1'b1;
17054: pixelout<=1'b1;
17055: pixelout<=1'b1;
17056: pixelout<=1'b1;
17057: pixelout<=1'b0;
17058: pixelout<=1'b0;
17059: pixelout<=1'b1;
17060: pixelout<=1'b1;
17061: pixelout<=1'b1;
17062: pixelout<=1'b1;
17063: pixelout<=1'b1;
17064: pixelout<=1'b1;
17065: pixelout<=1'b0;
17066: pixelout<=1'b0;
17067: pixelout<=1'b1;
17068: pixelout<=1'b1;
17069: pixelout<=1'b1;
17070: pixelout<=1'b1;
17071: pixelout<=1'b1;
17072: pixelout<=1'b1;
17073: pixelout<=1'b1;
17074: pixelout<=1'b1;
17075: pixelout<=1'b1;
17076: pixelout<=1'b1;
17077: pixelout<=1'b1;
17078: pixelout<=1'b1;
17079: pixelout<=1'b1;
17080: pixelout<=1'b1;
17081: pixelout<=1'b1;
17082: pixelout<=1'b1;
17083: pixelout<=1'b1;
17084: pixelout<=1'b1;
17085: pixelout<=1'b1;
17086: pixelout<=1'b1;
17087: pixelout<=1'b1;
17088: pixelout<=1'b1;
17089: pixelout<=1'b1;
17090: pixelout<=1'b1;
17091: pixelout<=1'b1;
17092: pixelout<=1'b1;
17093: pixelout<=1'b1;
17094: pixelout<=1'b1;
17095: pixelout<=1'b1;
17096: pixelout<=1'b1;
17097: pixelout<=1'b1;
17098: pixelout<=1'b1;
17099: pixelout<=1'b1;
17100: pixelout<=1'b1;
17101: pixelout<=1'b1;
17102: pixelout<=1'b1;
17103: pixelout<=1'b1;
17104: pixelout<=1'b1;
17105: pixelout<=1'b1;
17106: pixelout<=1'b1;
17107: pixelout<=1'b1;
17108: pixelout<=1'b1;
17109: pixelout<=1'b1;
17110: pixelout<=1'b1;
17111: pixelout<=1'b1;
17112: pixelout<=1'b0;
17113: pixelout<=1'b0;
17114: pixelout<=1'b1;
17115: pixelout<=1'b1;
17116: pixelout<=1'b1;
17117: pixelout<=1'b1;
17118: pixelout<=1'b0;
17119: pixelout<=1'b0;
17120: pixelout<=1'b1;
17121: pixelout<=1'b1;
17122: pixelout<=1'b1;
17123: pixelout<=1'b1;
17124: pixelout<=1'b1;
17125: pixelout<=1'b0;
17126: pixelout<=1'b0;
17127: pixelout<=1'b0;
17128: pixelout<=1'b0;
17129: pixelout<=1'b0;
17130: pixelout<=1'b1;
17131: pixelout<=1'b1;
17132: pixelout<=1'b1;
17133: pixelout<=1'b1;
17134: pixelout<=1'b1;
17135: pixelout<=1'b1;
17136: pixelout<=1'b1;
17137: pixelout<=1'b1;
17138: pixelout<=1'b1;
17139: pixelout<=1'b1;
17140: pixelout<=1'b1;
17141: pixelout<=1'b1;
17142: pixelout<=1'b1;
17143: pixelout<=1'b1;
17144: pixelout<=1'b1;
17145: pixelout<=1'b1;
17146: pixelout<=1'b1;
17147: pixelout<=1'b1;
17148: pixelout<=1'b1;
17149: pixelout<=1'b1;
17150: pixelout<=1'b1;
17151: pixelout<=1'b1;
17152: pixelout<=1'b1;
17153: pixelout<=1'b1;
17154: pixelout<=1'b1;
17155: pixelout<=1'b1;
17156: pixelout<=1'b1;
17157: pixelout<=1'b1;
17158: pixelout<=1'b1;
17159: pixelout<=1'b1;
17160: pixelout<=1'b1;
17161: pixelout<=1'b1;
17162: pixelout<=1'b1;
17163: pixelout<=1'b1;
17164: pixelout<=1'b1;
17165: pixelout<=1'b1;
17166: pixelout<=1'b1;
17167: pixelout<=1'b1;
17168: pixelout<=1'b1;
17169: pixelout<=1'b1;
17170: pixelout<=1'b1;
17171: pixelout<=1'b1;
17172: pixelout<=1'b1;
17173: pixelout<=1'b1;
17174: pixelout<=1'b1;
17175: pixelout<=1'b1;
17176: pixelout<=1'b1;
17177: pixelout<=1'b1;
17178: pixelout<=1'b1;
17179: pixelout<=1'b1;
17180: pixelout<=1'b1;
17181: pixelout<=1'b1;
17182: pixelout<=1'b1;
17183: pixelout<=1'b1;
17184: pixelout<=1'b1;
17185: pixelout<=1'b1;
17186: pixelout<=1'b1;
17187: pixelout<=1'b1;
17188: pixelout<=1'b1;
17189: pixelout<=1'b1;
17190: pixelout<=1'b1;
17191: pixelout<=1'b1;
17192: pixelout<=1'b1;
17193: pixelout<=1'b1;
17194: pixelout<=1'b1;
17195: pixelout<=1'b1;
17196: pixelout<=1'b1;
17197: pixelout<=1'b1;
17198: pixelout<=1'b1;
17199: pixelout<=1'b1;
17200: pixelout<=1'b1;
17201: pixelout<=1'b1;
17202: pixelout<=1'b1;
17203: pixelout<=1'b1;
17204: pixelout<=1'b1;
17205: pixelout<=1'b1;
17206: pixelout<=1'b1;
17207: pixelout<=1'b1;
17208: pixelout<=1'b1;
17209: pixelout<=1'b1;
17210: pixelout<=1'b1;
17211: pixelout<=1'b1;
17212: pixelout<=1'b1;
17213: pixelout<=1'b1;
17214: pixelout<=1'b1;
17215: pixelout<=1'b1;
17216: pixelout<=1'b1;
17217: pixelout<=1'b1;
17218: pixelout<=1'b1;
17219: pixelout<=1'b1;
17220: pixelout<=1'b1;
17221: pixelout<=1'b1;
17222: pixelout<=1'b1;
17223: pixelout<=1'b1;
17224: pixelout<=1'b0;
17225: pixelout<=1'b1;
17226: pixelout<=1'b1;
17227: pixelout<=1'b1;
17228: pixelout<=1'b1;
17229: pixelout<=1'b1;
17230: pixelout<=1'b1;
17231: pixelout<=1'b1;
17232: pixelout<=1'b1;
17233: pixelout<=1'b1;
17234: pixelout<=1'b1;
17235: pixelout<=1'b1;
17236: pixelout<=1'b1;
17237: pixelout<=1'b1;
17238: pixelout<=1'b1;
17239: pixelout<=1'b1;
17240: pixelout<=1'b1;
17241: pixelout<=1'b1;
17242: pixelout<=1'b1;
17243: pixelout<=1'b1;
17244: pixelout<=1'b1;
17245: pixelout<=1'b1;
17246: pixelout<=1'b1;
17247: pixelout<=1'b1;
17248: pixelout<=1'b1;
17249: pixelout<=1'b1;
17250: pixelout<=1'b1;
17251: pixelout<=1'b0;
17252: pixelout<=1'b0;
17253: pixelout<=1'b1;
17254: pixelout<=1'b1;
17255: pixelout<=1'b1;
17256: pixelout<=1'b1;
17257: pixelout<=1'b1;
17258: pixelout<=1'b1;
17259: pixelout<=1'b1;
17260: pixelout<=1'b1;
17261: pixelout<=1'b1;
17262: pixelout<=1'b1;
17263: pixelout<=1'b1;
17264: pixelout<=1'b1;
17265: pixelout<=1'b1;
17266: pixelout<=1'b1;
17267: pixelout<=1'b1;
17268: pixelout<=1'b1;
17269: pixelout<=1'b1;
17270: pixelout<=1'b1;
17271: pixelout<=1'b0;
17272: pixelout<=1'b1;
17273: pixelout<=1'b1;
17274: pixelout<=1'b1;
17275: pixelout<=1'b1;
17276: pixelout<=1'b1;
17277: pixelout<=1'b1;
17278: pixelout<=1'b1;
17279: pixelout<=1'b1;
17280: pixelout<=1'b1;
17281: pixelout<=1'b1;
17282: pixelout<=1'b1;
17283: pixelout<=1'b1;
17284: pixelout<=1'b1;
17285: pixelout<=1'b1;
17286: pixelout<=1'b1;
17287: pixelout<=1'b1;
17288: pixelout<=1'b1;
17289: pixelout<=1'b0;
17290: pixelout<=1'b1;
17291: pixelout<=1'b1;
17292: pixelout<=1'b1;
17293: pixelout<=1'b1;
17294: pixelout<=1'b1;
17295: pixelout<=1'b0;
17296: pixelout<=1'b1;
17297: pixelout<=1'b1;
17298: pixelout<=1'b1;
17299: pixelout<=1'b1;
17300: pixelout<=1'b1;
17301: pixelout<=1'b1;
17302: pixelout<=1'b1;
17303: pixelout<=1'b1;
17304: pixelout<=1'b1;
17305: pixelout<=1'b1;
17306: pixelout<=1'b1;
17307: pixelout<=1'b1;
17308: pixelout<=1'b0;
17309: pixelout<=1'b1;
17310: pixelout<=1'b1;
17311: pixelout<=1'b1;
17312: pixelout<=1'b1;
17313: pixelout<=1'b1;
17314: pixelout<=1'b1;
17315: pixelout<=1'b1;
17316: pixelout<=1'b1;
17317: pixelout<=1'b1;
17318: pixelout<=1'b1;
17319: pixelout<=1'b1;
17320: pixelout<=1'b1;
17321: pixelout<=1'b1;
17322: pixelout<=1'b1;
17323: pixelout<=1'b1;
17324: pixelout<=1'b1;
17325: pixelout<=1'b1;
17326: pixelout<=1'b1;
17327: pixelout<=1'b1;
17328: pixelout<=1'b1;
17329: pixelout<=1'b1;
17330: pixelout<=1'b1;
17331: pixelout<=1'b1;
17332: pixelout<=1'b1;
17333: pixelout<=1'b1;
17334: pixelout<=1'b1;
17335: pixelout<=1'b1;
17336: pixelout<=1'b1;
17337: pixelout<=1'b1;
17338: pixelout<=1'b1;
17339: pixelout<=1'b1;
17340: pixelout<=1'b1;
17341: pixelout<=1'b1;
17342: pixelout<=1'b1;
17343: pixelout<=1'b1;
17344: pixelout<=1'b1;
17345: pixelout<=1'b1;
17346: pixelout<=1'b1;
17347: pixelout<=1'b1;
17348: pixelout<=1'b1;
17349: pixelout<=1'b1;
17350: pixelout<=1'b0;
17351: pixelout<=1'b1;
17352: pixelout<=1'b1;
17353: pixelout<=1'b1;
17354: pixelout<=1'b1;
17355: pixelout<=1'b1;
17356: pixelout<=1'b1;
17357: pixelout<=1'b1;
17358: pixelout<=1'b1;
17359: pixelout<=1'b1;
17360: pixelout<=1'b1;
17361: pixelout<=1'b0;
17362: pixelout<=1'b1;
17363: pixelout<=1'b1;
17364: pixelout<=1'b1;
17365: pixelout<=1'b1;
17366: pixelout<=1'b1;
17367: pixelout<=1'b0;
17368: pixelout<=1'b1;
17369: pixelout<=1'b1;
17370: pixelout<=1'b1;
17371: pixelout<=1'b1;
17372: pixelout<=1'b1;
17373: pixelout<=1'b1;
17374: pixelout<=1'b1;
17375: pixelout<=1'b1;
17376: pixelout<=1'b1;
17377: pixelout<=1'b1;
17378: pixelout<=1'b1;
17379: pixelout<=1'b1;
17380: pixelout<=1'b1;
17381: pixelout<=1'b1;
17382: pixelout<=1'b1;
17383: pixelout<=1'b1;
17384: pixelout<=1'b1;
17385: pixelout<=1'b1;
17386: pixelout<=1'b1;
17387: pixelout<=1'b1;
17388: pixelout<=1'b1;
17389: pixelout<=1'b1;
17390: pixelout<=1'b1;
17391: pixelout<=1'b1;
17392: pixelout<=1'b1;
17393: pixelout<=1'b1;
17394: pixelout<=1'b1;
17395: pixelout<=1'b1;
17396: pixelout<=1'b1;
17397: pixelout<=1'b1;
17398: pixelout<=1'b1;
17399: pixelout<=1'b1;
17400: pixelout<=1'b1;
17401: pixelout<=1'b1;
17402: pixelout<=1'b1;
17403: pixelout<=1'b1;
17404: pixelout<=1'b1;
17405: pixelout<=1'b1;
17406: pixelout<=1'b1;
17407: pixelout<=1'b1;
17408: pixelout<=1'b1;
17409: pixelout<=1'b1;
17410: pixelout<=1'b1;
17411: pixelout<=1'b1;
17412: pixelout<=1'b1;
17413: pixelout<=1'b1;
17414: pixelout<=1'b1;
17415: pixelout<=1'b1;
17416: pixelout<=1'b1;
17417: pixelout<=1'b1;
17418: pixelout<=1'b1;
17419: pixelout<=1'b1;
17420: pixelout<=1'b1;
17421: pixelout<=1'b1;
17422: pixelout<=1'b1;
17423: pixelout<=1'b1;
17424: pixelout<=1'b1;
17425: pixelout<=1'b1;
17426: pixelout<=1'b1;
17427: pixelout<=1'b1;
17428: pixelout<=1'b1;
17429: pixelout<=1'b1;
17430: pixelout<=1'b1;
17431: pixelout<=1'b1;
17432: pixelout<=1'b1;
17433: pixelout<=1'b1;
17434: pixelout<=1'b1;
17435: pixelout<=1'b1;
17436: pixelout<=1'b1;
17437: pixelout<=1'b1;
17438: pixelout<=1'b1;
17439: pixelout<=1'b1;
17440: pixelout<=1'b1;
17441: pixelout<=1'b1;
17442: pixelout<=1'b1;
17443: pixelout<=1'b1;
17444: pixelout<=1'b1;
17445: pixelout<=1'b1;
17446: pixelout<=1'b1;
17447: pixelout<=1'b1;
17448: pixelout<=1'b1;
17449: pixelout<=1'b1;
17450: pixelout<=1'b1;
17451: pixelout<=1'b1;
17452: pixelout<=1'b1;
17453: pixelout<=1'b1;
17454: pixelout<=1'b1;
17455: pixelout<=1'b1;
17456: pixelout<=1'b1;
17457: pixelout<=1'b1;
17458: pixelout<=1'b1;
17459: pixelout<=1'b1;
17460: pixelout<=1'b1;
17461: pixelout<=1'b1;
17462: pixelout<=1'b1;
17463: pixelout<=1'b1;
17464: pixelout<=1'b0;
17465: pixelout<=1'b1;
17466: pixelout<=1'b1;
17467: pixelout<=1'b1;
17468: pixelout<=1'b1;
17469: pixelout<=1'b1;
17470: pixelout<=1'b1;
17471: pixelout<=1'b1;
17472: pixelout<=1'b1;
17473: pixelout<=1'b1;
17474: pixelout<=1'b1;
17475: pixelout<=1'b1;
17476: pixelout<=1'b1;
17477: pixelout<=1'b1;
17478: pixelout<=1'b1;
17479: pixelout<=1'b1;
17480: pixelout<=1'b1;
17481: pixelout<=1'b1;
17482: pixelout<=1'b1;
17483: pixelout<=1'b1;
17484: pixelout<=1'b1;
17485: pixelout<=1'b1;
17486: pixelout<=1'b1;
17487: pixelout<=1'b1;
17488: pixelout<=1'b1;
17489: pixelout<=1'b1;
17490: pixelout<=1'b1;
17491: pixelout<=1'b1;
17492: pixelout<=1'b0;
17493: pixelout<=1'b1;
17494: pixelout<=1'b1;
17495: pixelout<=1'b1;
17496: pixelout<=1'b1;
17497: pixelout<=1'b1;
17498: pixelout<=1'b1;
17499: pixelout<=1'b1;
17500: pixelout<=1'b1;
17501: pixelout<=1'b1;
17502: pixelout<=1'b1;
17503: pixelout<=1'b1;
17504: pixelout<=1'b1;
17505: pixelout<=1'b1;
17506: pixelout<=1'b1;
17507: pixelout<=1'b1;
17508: pixelout<=1'b1;
17509: pixelout<=1'b1;
17510: pixelout<=1'b1;
17511: pixelout<=1'b0;
17512: pixelout<=1'b1;
17513: pixelout<=1'b1;
17514: pixelout<=1'b1;
17515: pixelout<=1'b1;
17516: pixelout<=1'b1;
17517: pixelout<=1'b1;
17518: pixelout<=1'b1;
17519: pixelout<=1'b1;
17520: pixelout<=1'b1;
17521: pixelout<=1'b1;
17522: pixelout<=1'b1;
17523: pixelout<=1'b1;
17524: pixelout<=1'b1;
17525: pixelout<=1'b1;
17526: pixelout<=1'b1;
17527: pixelout<=1'b1;
17528: pixelout<=1'b1;
17529: pixelout<=1'b0;
17530: pixelout<=1'b1;
17531: pixelout<=1'b1;
17532: pixelout<=1'b1;
17533: pixelout<=1'b1;
17534: pixelout<=1'b1;
17535: pixelout<=1'b0;
17536: pixelout<=1'b1;
17537: pixelout<=1'b1;
17538: pixelout<=1'b1;
17539: pixelout<=1'b1;
17540: pixelout<=1'b1;
17541: pixelout<=1'b1;
17542: pixelout<=1'b1;
17543: pixelout<=1'b1;
17544: pixelout<=1'b1;
17545: pixelout<=1'b1;
17546: pixelout<=1'b1;
17547: pixelout<=1'b1;
17548: pixelout<=1'b0;
17549: pixelout<=1'b1;
17550: pixelout<=1'b1;
17551: pixelout<=1'b1;
17552: pixelout<=1'b1;
17553: pixelout<=1'b1;
17554: pixelout<=1'b1;
17555: pixelout<=1'b1;
17556: pixelout<=1'b1;
17557: pixelout<=1'b1;
17558: pixelout<=1'b1;
17559: pixelout<=1'b1;
17560: pixelout<=1'b1;
17561: pixelout<=1'b1;
17562: pixelout<=1'b1;
17563: pixelout<=1'b1;
17564: pixelout<=1'b1;
17565: pixelout<=1'b1;
17566: pixelout<=1'b1;
17567: pixelout<=1'b1;
17568: pixelout<=1'b1;
17569: pixelout<=1'b1;
17570: pixelout<=1'b1;
17571: pixelout<=1'b1;
17572: pixelout<=1'b1;
17573: pixelout<=1'b1;
17574: pixelout<=1'b1;
17575: pixelout<=1'b1;
17576: pixelout<=1'b1;
17577: pixelout<=1'b1;
17578: pixelout<=1'b1;
17579: pixelout<=1'b1;
17580: pixelout<=1'b1;
17581: pixelout<=1'b1;
17582: pixelout<=1'b1;
17583: pixelout<=1'b1;
17584: pixelout<=1'b1;
17585: pixelout<=1'b1;
17586: pixelout<=1'b1;
17587: pixelout<=1'b1;
17588: pixelout<=1'b1;
17589: pixelout<=1'b1;
17590: pixelout<=1'b0;
17591: pixelout<=1'b1;
17592: pixelout<=1'b1;
17593: pixelout<=1'b1;
17594: pixelout<=1'b1;
17595: pixelout<=1'b1;
17596: pixelout<=1'b1;
17597: pixelout<=1'b1;
17598: pixelout<=1'b1;
17599: pixelout<=1'b1;
17600: pixelout<=1'b1;
17601: pixelout<=1'b0;
17602: pixelout<=1'b1;
17603: pixelout<=1'b1;
17604: pixelout<=1'b1;
17605: pixelout<=1'b1;
17606: pixelout<=1'b1;
17607: pixelout<=1'b0;
17608: pixelout<=1'b1;
17609: pixelout<=1'b1;
17610: pixelout<=1'b1;
17611: pixelout<=1'b1;
17612: pixelout<=1'b1;
17613: pixelout<=1'b1;
17614: pixelout<=1'b1;
17615: pixelout<=1'b1;
17616: pixelout<=1'b1;
17617: pixelout<=1'b1;
17618: pixelout<=1'b1;
17619: pixelout<=1'b1;
17620: pixelout<=1'b1;
17621: pixelout<=1'b1;
17622: pixelout<=1'b1;
17623: pixelout<=1'b1;
17624: pixelout<=1'b1;
17625: pixelout<=1'b1;
17626: pixelout<=1'b1;
17627: pixelout<=1'b1;
17628: pixelout<=1'b1;
17629: pixelout<=1'b1;
17630: pixelout<=1'b1;
17631: pixelout<=1'b1;
17632: pixelout<=1'b1;
17633: pixelout<=1'b1;
17634: pixelout<=1'b1;
17635: pixelout<=1'b1;
17636: pixelout<=1'b1;
17637: pixelout<=1'b1;
17638: pixelout<=1'b1;
17639: pixelout<=1'b1;
17640: pixelout<=1'b1;
17641: pixelout<=1'b1;
17642: pixelout<=1'b1;
17643: pixelout<=1'b1;
17644: pixelout<=1'b1;
17645: pixelout<=1'b1;
17646: pixelout<=1'b1;
17647: pixelout<=1'b1;
17648: pixelout<=1'b1;
17649: pixelout<=1'b1;
17650: pixelout<=1'b1;
17651: pixelout<=1'b1;
17652: pixelout<=1'b1;
17653: pixelout<=1'b1;
17654: pixelout<=1'b1;
17655: pixelout<=1'b1;
17656: pixelout<=1'b1;
17657: pixelout<=1'b1;
17658: pixelout<=1'b1;
17659: pixelout<=1'b1;
17660: pixelout<=1'b1;
17661: pixelout<=1'b1;
17662: pixelout<=1'b1;
17663: pixelout<=1'b1;
17664: pixelout<=1'b1;
17665: pixelout<=1'b1;
17666: pixelout<=1'b1;
17667: pixelout<=1'b1;
17668: pixelout<=1'b1;
17669: pixelout<=1'b1;
17670: pixelout<=1'b1;
17671: pixelout<=1'b1;
17672: pixelout<=1'b1;
17673: pixelout<=1'b1;
17674: pixelout<=1'b1;
17675: pixelout<=1'b1;
17676: pixelout<=1'b1;
17677: pixelout<=1'b1;
17678: pixelout<=1'b1;
17679: pixelout<=1'b1;
17680: pixelout<=1'b1;
17681: pixelout<=1'b1;
17682: pixelout<=1'b1;
17683: pixelout<=1'b1;
17684: pixelout<=1'b1;
17685: pixelout<=1'b1;
17686: pixelout<=1'b1;
17687: pixelout<=1'b1;
17688: pixelout<=1'b1;
17689: pixelout<=1'b1;
17690: pixelout<=1'b1;
17691: pixelout<=1'b1;
17692: pixelout<=1'b1;
17693: pixelout<=1'b1;
17694: pixelout<=1'b1;
17695: pixelout<=1'b1;
17696: pixelout<=1'b1;
17697: pixelout<=1'b1;
17698: pixelout<=1'b1;
17699: pixelout<=1'b1;
17700: pixelout<=1'b1;
17701: pixelout<=1'b1;
17702: pixelout<=1'b1;
17703: pixelout<=1'b1;
17704: pixelout<=1'b0;
17705: pixelout<=1'b1;
17706: pixelout<=1'b1;
17707: pixelout<=1'b1;
17708: pixelout<=1'b1;
17709: pixelout<=1'b1;
17710: pixelout<=1'b1;
17711: pixelout<=1'b1;
17712: pixelout<=1'b1;
17713: pixelout<=1'b1;
17714: pixelout<=1'b1;
17715: pixelout<=1'b1;
17716: pixelout<=1'b1;
17717: pixelout<=1'b1;
17718: pixelout<=1'b1;
17719: pixelout<=1'b1;
17720: pixelout<=1'b1;
17721: pixelout<=1'b1;
17722: pixelout<=1'b1;
17723: pixelout<=1'b1;
17724: pixelout<=1'b1;
17725: pixelout<=1'b1;
17726: pixelout<=1'b1;
17727: pixelout<=1'b1;
17728: pixelout<=1'b1;
17729: pixelout<=1'b1;
17730: pixelout<=1'b1;
17731: pixelout<=1'b1;
17732: pixelout<=1'b0;
17733: pixelout<=1'b1;
17734: pixelout<=1'b1;
17735: pixelout<=1'b1;
17736: pixelout<=1'b1;
17737: pixelout<=1'b1;
17738: pixelout<=1'b1;
17739: pixelout<=1'b1;
17740: pixelout<=1'b1;
17741: pixelout<=1'b1;
17742: pixelout<=1'b1;
17743: pixelout<=1'b1;
17744: pixelout<=1'b1;
17745: pixelout<=1'b1;
17746: pixelout<=1'b1;
17747: pixelout<=1'b1;
17748: pixelout<=1'b1;
17749: pixelout<=1'b1;
17750: pixelout<=1'b1;
17751: pixelout<=1'b0;
17752: pixelout<=1'b1;
17753: pixelout<=1'b1;
17754: pixelout<=1'b1;
17755: pixelout<=1'b1;
17756: pixelout<=1'b1;
17757: pixelout<=1'b1;
17758: pixelout<=1'b1;
17759: pixelout<=1'b1;
17760: pixelout<=1'b1;
17761: pixelout<=1'b1;
17762: pixelout<=1'b1;
17763: pixelout<=1'b1;
17764: pixelout<=1'b1;
17765: pixelout<=1'b1;
17766: pixelout<=1'b1;
17767: pixelout<=1'b1;
17768: pixelout<=1'b1;
17769: pixelout<=1'b0;
17770: pixelout<=1'b1;
17771: pixelout<=1'b1;
17772: pixelout<=1'b1;
17773: pixelout<=1'b1;
17774: pixelout<=1'b1;
17775: pixelout<=1'b0;
17776: pixelout<=1'b1;
17777: pixelout<=1'b1;
17778: pixelout<=1'b1;
17779: pixelout<=1'b1;
17780: pixelout<=1'b1;
17781: pixelout<=1'b1;
17782: pixelout<=1'b1;
17783: pixelout<=1'b1;
17784: pixelout<=1'b1;
17785: pixelout<=1'b1;
17786: pixelout<=1'b1;
17787: pixelout<=1'b1;
17788: pixelout<=1'b0;
17789: pixelout<=1'b1;
17790: pixelout<=1'b0;
17791: pixelout<=1'b0;
17792: pixelout<=1'b0;
17793: pixelout<=1'b1;
17794: pixelout<=1'b1;
17795: pixelout<=1'b0;
17796: pixelout<=1'b1;
17797: pixelout<=1'b1;
17798: pixelout<=1'b0;
17799: pixelout<=1'b1;
17800: pixelout<=1'b1;
17801: pixelout<=1'b0;
17802: pixelout<=1'b0;
17803: pixelout<=1'b0;
17804: pixelout<=1'b0;
17805: pixelout<=1'b1;
17806: pixelout<=1'b1;
17807: pixelout<=1'b0;
17808: pixelout<=1'b0;
17809: pixelout<=1'b0;
17810: pixelout<=1'b1;
17811: pixelout<=1'b1;
17812: pixelout<=1'b1;
17813: pixelout<=1'b0;
17814: pixelout<=1'b1;
17815: pixelout<=1'b1;
17816: pixelout<=1'b1;
17817: pixelout<=1'b0;
17818: pixelout<=1'b1;
17819: pixelout<=1'b1;
17820: pixelout<=1'b0;
17821: pixelout<=1'b0;
17822: pixelout<=1'b0;
17823: pixelout<=1'b0;
17824: pixelout<=1'b1;
17825: pixelout<=1'b1;
17826: pixelout<=1'b1;
17827: pixelout<=1'b1;
17828: pixelout<=1'b1;
17829: pixelout<=1'b1;
17830: pixelout<=1'b0;
17831: pixelout<=1'b1;
17832: pixelout<=1'b1;
17833: pixelout<=1'b1;
17834: pixelout<=1'b1;
17835: pixelout<=1'b1;
17836: pixelout<=1'b1;
17837: pixelout<=1'b1;
17838: pixelout<=1'b1;
17839: pixelout<=1'b1;
17840: pixelout<=1'b1;
17841: pixelout<=1'b0;
17842: pixelout<=1'b1;
17843: pixelout<=1'b1;
17844: pixelout<=1'b1;
17845: pixelout<=1'b1;
17846: pixelout<=1'b1;
17847: pixelout<=1'b0;
17848: pixelout<=1'b1;
17849: pixelout<=1'b1;
17850: pixelout<=1'b1;
17851: pixelout<=1'b1;
17852: pixelout<=1'b1;
17853: pixelout<=1'b0;
17854: pixelout<=1'b0;
17855: pixelout<=1'b0;
17856: pixelout<=1'b1;
17857: pixelout<=1'b1;
17858: pixelout<=1'b0;
17859: pixelout<=1'b0;
17860: pixelout<=1'b1;
17861: pixelout<=1'b1;
17862: pixelout<=1'b1;
17863: pixelout<=1'b1;
17864: pixelout<=1'b1;
17865: pixelout<=1'b1;
17866: pixelout<=1'b1;
17867: pixelout<=1'b1;
17868: pixelout<=1'b1;
17869: pixelout<=1'b0;
17870: pixelout<=1'b0;
17871: pixelout<=1'b0;
17872: pixelout<=1'b0;
17873: pixelout<=1'b1;
17874: pixelout<=1'b0;
17875: pixelout<=1'b0;
17876: pixelout<=1'b0;
17877: pixelout<=1'b1;
17878: pixelout<=1'b1;
17879: pixelout<=1'b1;
17880: pixelout<=1'b1;
17881: pixelout<=1'b0;
17882: pixelout<=1'b0;
17883: pixelout<=1'b0;
17884: pixelout<=1'b1;
17885: pixelout<=1'b1;
17886: pixelout<=1'b1;
17887: pixelout<=1'b1;
17888: pixelout<=1'b1;
17889: pixelout<=1'b0;
17890: pixelout<=1'b0;
17891: pixelout<=1'b0;
17892: pixelout<=1'b1;
17893: pixelout<=1'b1;
17894: pixelout<=1'b0;
17895: pixelout<=1'b1;
17896: pixelout<=1'b1;
17897: pixelout<=1'b1;
17898: pixelout<=1'b0;
17899: pixelout<=1'b1;
17900: pixelout<=1'b1;
17901: pixelout<=1'b1;
17902: pixelout<=1'b0;
17903: pixelout<=1'b0;
17904: pixelout<=1'b1;
17905: pixelout<=1'b1;
17906: pixelout<=1'b1;
17907: pixelout<=1'b1;
17908: pixelout<=1'b1;
17909: pixelout<=1'b0;
17910: pixelout<=1'b1;
17911: pixelout<=1'b1;
17912: pixelout<=1'b1;
17913: pixelout<=1'b1;
17914: pixelout<=1'b1;
17915: pixelout<=1'b1;
17916: pixelout<=1'b0;
17917: pixelout<=1'b1;
17918: pixelout<=1'b1;
17919: pixelout<=1'b0;
17920: pixelout<=1'b0;
17921: pixelout<=1'b0;
17922: pixelout<=1'b1;
17923: pixelout<=1'b1;
17924: pixelout<=1'b0;
17925: pixelout<=1'b0;
17926: pixelout<=1'b0;
17927: pixelout<=1'b1;
17928: pixelout<=1'b1;
17929: pixelout<=1'b1;
17930: pixelout<=1'b1;
17931: pixelout<=1'b0;
17932: pixelout<=1'b0;
17933: pixelout<=1'b1;
17934: pixelout<=1'b1;
17935: pixelout<=1'b1;
17936: pixelout<=1'b1;
17937: pixelout<=1'b1;
17938: pixelout<=1'b0;
17939: pixelout<=1'b1;
17940: pixelout<=1'b0;
17941: pixelout<=1'b1;
17942: pixelout<=1'b0;
17943: pixelout<=1'b1;
17944: pixelout<=1'b0;
17945: pixelout<=1'b0;
17946: pixelout<=1'b0;
17947: pixelout<=1'b0;
17948: pixelout<=1'b1;
17949: pixelout<=1'b1;
17950: pixelout<=1'b1;
17951: pixelout<=1'b1;
17952: pixelout<=1'b0;
17953: pixelout<=1'b0;
17954: pixelout<=1'b1;
17955: pixelout<=1'b1;
17956: pixelout<=1'b1;
17957: pixelout<=1'b1;
17958: pixelout<=1'b1;
17959: pixelout<=1'b0;
17960: pixelout<=1'b0;
17961: pixelout<=1'b0;
17962: pixelout<=1'b1;
17963: pixelout<=1'b1;
17964: pixelout<=1'b1;
17965: pixelout<=1'b1;
17966: pixelout<=1'b0;
17967: pixelout<=1'b0;
17968: pixelout<=1'b0;
17969: pixelout<=1'b1;
17970: pixelout<=1'b1;
17971: pixelout<=1'b1;
17972: pixelout<=1'b0;
17973: pixelout<=1'b1;
17974: pixelout<=1'b0;
17975: pixelout<=1'b0;
17976: pixelout<=1'b0;
17977: pixelout<=1'b0;
17978: pixelout<=1'b1;
17979: pixelout<=1'b1;
17980: pixelout<=1'b1;
17981: pixelout<=1'b1;
17982: pixelout<=1'b0;
17983: pixelout<=1'b0;
17984: pixelout<=1'b1;
17985: pixelout<=1'b1;
17986: pixelout<=1'b1;
17987: pixelout<=1'b1;
17988: pixelout<=1'b0;
17989: pixelout<=1'b0;
17990: pixelout<=1'b0;
17991: pixelout<=1'b0;
17992: pixelout<=1'b1;
17993: pixelout<=1'b1;
17994: pixelout<=1'b1;
17995: pixelout<=1'b1;
17996: pixelout<=1'b1;
17997: pixelout<=1'b1;
17998: pixelout<=1'b1;
17999: pixelout<=1'b1;
18000: pixelout<=1'b1;
18001: pixelout<=1'b1;
18002: pixelout<=1'b1;
18003: pixelout<=1'b1;
18004: pixelout<=1'b1;
18005: pixelout<=1'b1;
18006: pixelout<=1'b1;
18007: pixelout<=1'b1;
18008: pixelout<=1'b1;
18009: pixelout<=1'b0;
18010: pixelout<=1'b1;
18011: pixelout<=1'b1;
18012: pixelout<=1'b1;
18013: pixelout<=1'b1;
18014: pixelout<=1'b1;
18015: pixelout<=1'b0;
18016: pixelout<=1'b0;
18017: pixelout<=1'b0;
18018: pixelout<=1'b0;
18019: pixelout<=1'b0;
18020: pixelout<=1'b1;
18021: pixelout<=1'b1;
18022: pixelout<=1'b1;
18023: pixelout<=1'b1;
18024: pixelout<=1'b0;
18025: pixelout<=1'b0;
18026: pixelout<=1'b0;
18027: pixelout<=1'b0;
18028: pixelout<=1'b0;
18029: pixelout<=1'b1;
18030: pixelout<=1'b0;
18031: pixelout<=1'b1;
18032: pixelout<=1'b1;
18033: pixelout<=1'b0;
18034: pixelout<=1'b1;
18035: pixelout<=1'b0;
18036: pixelout<=1'b1;
18037: pixelout<=1'b1;
18038: pixelout<=1'b0;
18039: pixelout<=1'b1;
18040: pixelout<=1'b1;
18041: pixelout<=1'b0;
18042: pixelout<=1'b1;
18043: pixelout<=1'b1;
18044: pixelout<=1'b1;
18045: pixelout<=1'b1;
18046: pixelout<=1'b1;
18047: pixelout<=1'b1;
18048: pixelout<=1'b1;
18049: pixelout<=1'b1;
18050: pixelout<=1'b1;
18051: pixelout<=1'b0;
18052: pixelout<=1'b1;
18053: pixelout<=1'b0;
18054: pixelout<=1'b1;
18055: pixelout<=1'b1;
18056: pixelout<=1'b1;
18057: pixelout<=1'b0;
18058: pixelout<=1'b1;
18059: pixelout<=1'b0;
18060: pixelout<=1'b1;
18061: pixelout<=1'b1;
18062: pixelout<=1'b1;
18063: pixelout<=1'b0;
18064: pixelout<=1'b1;
18065: pixelout<=1'b1;
18066: pixelout<=1'b1;
18067: pixelout<=1'b1;
18068: pixelout<=1'b1;
18069: pixelout<=1'b1;
18070: pixelout<=1'b0;
18071: pixelout<=1'b1;
18072: pixelout<=1'b1;
18073: pixelout<=1'b1;
18074: pixelout<=1'b1;
18075: pixelout<=1'b1;
18076: pixelout<=1'b1;
18077: pixelout<=1'b0;
18078: pixelout<=1'b0;
18079: pixelout<=1'b0;
18080: pixelout<=1'b0;
18081: pixelout<=1'b0;
18082: pixelout<=1'b1;
18083: pixelout<=1'b1;
18084: pixelout<=1'b1;
18085: pixelout<=1'b1;
18086: pixelout<=1'b1;
18087: pixelout<=1'b0;
18088: pixelout<=1'b1;
18089: pixelout<=1'b1;
18090: pixelout<=1'b1;
18091: pixelout<=1'b0;
18092: pixelout<=1'b1;
18093: pixelout<=1'b1;
18094: pixelout<=1'b1;
18095: pixelout<=1'b1;
18096: pixelout<=1'b1;
18097: pixelout<=1'b1;
18098: pixelout<=1'b1;
18099: pixelout<=1'b1;
18100: pixelout<=1'b1;
18101: pixelout<=1'b0;
18102: pixelout<=1'b1;
18103: pixelout<=1'b1;
18104: pixelout<=1'b1;
18105: pixelout<=1'b1;
18106: pixelout<=1'b1;
18107: pixelout<=1'b1;
18108: pixelout<=1'b0;
18109: pixelout<=1'b1;
18110: pixelout<=1'b1;
18111: pixelout<=1'b1;
18112: pixelout<=1'b0;
18113: pixelout<=1'b1;
18114: pixelout<=1'b0;
18115: pixelout<=1'b1;
18116: pixelout<=1'b1;
18117: pixelout<=1'b0;
18118: pixelout<=1'b1;
18119: pixelout<=1'b0;
18120: pixelout<=1'b1;
18121: pixelout<=1'b1;
18122: pixelout<=1'b1;
18123: pixelout<=1'b1;
18124: pixelout<=1'b1;
18125: pixelout<=1'b1;
18126: pixelout<=1'b1;
18127: pixelout<=1'b1;
18128: pixelout<=1'b0;
18129: pixelout<=1'b1;
18130: pixelout<=1'b1;
18131: pixelout<=1'b1;
18132: pixelout<=1'b0;
18133: pixelout<=1'b1;
18134: pixelout<=1'b0;
18135: pixelout<=1'b1;
18136: pixelout<=1'b1;
18137: pixelout<=1'b1;
18138: pixelout<=1'b0;
18139: pixelout<=1'b1;
18140: pixelout<=1'b0;
18141: pixelout<=1'b1;
18142: pixelout<=1'b1;
18143: pixelout<=1'b1;
18144: pixelout<=1'b1;
18145: pixelout<=1'b1;
18146: pixelout<=1'b1;
18147: pixelout<=1'b0;
18148: pixelout<=1'b1;
18149: pixelout<=1'b1;
18150: pixelout<=1'b1;
18151: pixelout<=1'b1;
18152: pixelout<=1'b1;
18153: pixelout<=1'b1;
18154: pixelout<=1'b1;
18155: pixelout<=1'b1;
18156: pixelout<=1'b0;
18157: pixelout<=1'b1;
18158: pixelout<=1'b0;
18159: pixelout<=1'b1;
18160: pixelout<=1'b1;
18161: pixelout<=1'b1;
18162: pixelout<=1'b0;
18163: pixelout<=1'b1;
18164: pixelout<=1'b0;
18165: pixelout<=1'b1;
18166: pixelout<=1'b1;
18167: pixelout<=1'b0;
18168: pixelout<=1'b1;
18169: pixelout<=1'b0;
18170: pixelout<=1'b1;
18171: pixelout<=1'b1;
18172: pixelout<=1'b1;
18173: pixelout<=1'b1;
18174: pixelout<=1'b1;
18175: pixelout<=1'b1;
18176: pixelout<=1'b1;
18177: pixelout<=1'b1;
18178: pixelout<=1'b0;
18179: pixelout<=1'b1;
18180: pixelout<=1'b0;
18181: pixelout<=1'b1;
18182: pixelout<=1'b0;
18183: pixelout<=1'b1;
18184: pixelout<=1'b0;
18185: pixelout<=1'b1;
18186: pixelout<=1'b1;
18187: pixelout<=1'b1;
18188: pixelout<=1'b0;
18189: pixelout<=1'b1;
18190: pixelout<=1'b0;
18191: pixelout<=1'b1;
18192: pixelout<=1'b1;
18193: pixelout<=1'b1;
18194: pixelout<=1'b1;
18195: pixelout<=1'b1;
18196: pixelout<=1'b1;
18197: pixelout<=1'b1;
18198: pixelout<=1'b1;
18199: pixelout<=1'b1;
18200: pixelout<=1'b1;
18201: pixelout<=1'b1;
18202: pixelout<=1'b1;
18203: pixelout<=1'b0;
18204: pixelout<=1'b1;
18205: pixelout<=1'b0;
18206: pixelout<=1'b1;
18207: pixelout<=1'b1;
18208: pixelout<=1'b1;
18209: pixelout<=1'b0;
18210: pixelout<=1'b1;
18211: pixelout<=1'b1;
18212: pixelout<=1'b0;
18213: pixelout<=1'b1;
18214: pixelout<=1'b0;
18215: pixelout<=1'b1;
18216: pixelout<=1'b1;
18217: pixelout<=1'b1;
18218: pixelout<=1'b0;
18219: pixelout<=1'b1;
18220: pixelout<=1'b0;
18221: pixelout<=1'b1;
18222: pixelout<=1'b1;
18223: pixelout<=1'b1;
18224: pixelout<=1'b1;
18225: pixelout<=1'b1;
18226: pixelout<=1'b1;
18227: pixelout<=1'b1;
18228: pixelout<=1'b1;
18229: pixelout<=1'b1;
18230: pixelout<=1'b1;
18231: pixelout<=1'b0;
18232: pixelout<=1'b1;
18233: pixelout<=1'b1;
18234: pixelout<=1'b1;
18235: pixelout<=1'b1;
18236: pixelout<=1'b1;
18237: pixelout<=1'b1;
18238: pixelout<=1'b1;
18239: pixelout<=1'b1;
18240: pixelout<=1'b1;
18241: pixelout<=1'b1;
18242: pixelout<=1'b1;
18243: pixelout<=1'b1;
18244: pixelout<=1'b1;
18245: pixelout<=1'b1;
18246: pixelout<=1'b1;
18247: pixelout<=1'b1;
18248: pixelout<=1'b1;
18249: pixelout<=1'b0;
18250: pixelout<=1'b1;
18251: pixelout<=1'b1;
18252: pixelout<=1'b1;
18253: pixelout<=1'b1;
18254: pixelout<=1'b1;
18255: pixelout<=1'b0;
18256: pixelout<=1'b1;
18257: pixelout<=1'b1;
18258: pixelout<=1'b1;
18259: pixelout<=1'b1;
18260: pixelout<=1'b1;
18261: pixelout<=1'b1;
18262: pixelout<=1'b1;
18263: pixelout<=1'b1;
18264: pixelout<=1'b1;
18265: pixelout<=1'b1;
18266: pixelout<=1'b1;
18267: pixelout<=1'b1;
18268: pixelout<=1'b0;
18269: pixelout<=1'b1;
18270: pixelout<=1'b0;
18271: pixelout<=1'b1;
18272: pixelout<=1'b1;
18273: pixelout<=1'b0;
18274: pixelout<=1'b1;
18275: pixelout<=1'b0;
18276: pixelout<=1'b1;
18277: pixelout<=1'b1;
18278: pixelout<=1'b0;
18279: pixelout<=1'b1;
18280: pixelout<=1'b1;
18281: pixelout<=1'b1;
18282: pixelout<=1'b0;
18283: pixelout<=1'b0;
18284: pixelout<=1'b1;
18285: pixelout<=1'b1;
18286: pixelout<=1'b1;
18287: pixelout<=1'b1;
18288: pixelout<=1'b1;
18289: pixelout<=1'b1;
18290: pixelout<=1'b1;
18291: pixelout<=1'b0;
18292: pixelout<=1'b1;
18293: pixelout<=1'b0;
18294: pixelout<=1'b1;
18295: pixelout<=1'b1;
18296: pixelout<=1'b1;
18297: pixelout<=1'b0;
18298: pixelout<=1'b1;
18299: pixelout<=1'b0;
18300: pixelout<=1'b1;
18301: pixelout<=1'b1;
18302: pixelout<=1'b1;
18303: pixelout<=1'b0;
18304: pixelout<=1'b1;
18305: pixelout<=1'b1;
18306: pixelout<=1'b1;
18307: pixelout<=1'b1;
18308: pixelout<=1'b1;
18309: pixelout<=1'b1;
18310: pixelout<=1'b0;
18311: pixelout<=1'b1;
18312: pixelout<=1'b1;
18313: pixelout<=1'b1;
18314: pixelout<=1'b1;
18315: pixelout<=1'b1;
18316: pixelout<=1'b1;
18317: pixelout<=1'b1;
18318: pixelout<=1'b1;
18319: pixelout<=1'b1;
18320: pixelout<=1'b1;
18321: pixelout<=1'b0;
18322: pixelout<=1'b1;
18323: pixelout<=1'b1;
18324: pixelout<=1'b1;
18325: pixelout<=1'b1;
18326: pixelout<=1'b1;
18327: pixelout<=1'b0;
18328: pixelout<=1'b1;
18329: pixelout<=1'b1;
18330: pixelout<=1'b1;
18331: pixelout<=1'b0;
18332: pixelout<=1'b1;
18333: pixelout<=1'b1;
18334: pixelout<=1'b1;
18335: pixelout<=1'b1;
18336: pixelout<=1'b1;
18337: pixelout<=1'b1;
18338: pixelout<=1'b1;
18339: pixelout<=1'b1;
18340: pixelout<=1'b1;
18341: pixelout<=1'b0;
18342: pixelout<=1'b1;
18343: pixelout<=1'b1;
18344: pixelout<=1'b1;
18345: pixelout<=1'b1;
18346: pixelout<=1'b1;
18347: pixelout<=1'b1;
18348: pixelout<=1'b0;
18349: pixelout<=1'b1;
18350: pixelout<=1'b1;
18351: pixelout<=1'b1;
18352: pixelout<=1'b0;
18353: pixelout<=1'b1;
18354: pixelout<=1'b0;
18355: pixelout<=1'b1;
18356: pixelout<=1'b1;
18357: pixelout<=1'b0;
18358: pixelout<=1'b1;
18359: pixelout<=1'b0;
18360: pixelout<=1'b1;
18361: pixelout<=1'b1;
18362: pixelout<=1'b1;
18363: pixelout<=1'b1;
18364: pixelout<=1'b1;
18365: pixelout<=1'b1;
18366: pixelout<=1'b1;
18367: pixelout<=1'b1;
18368: pixelout<=1'b0;
18369: pixelout<=1'b0;
18370: pixelout<=1'b0;
18371: pixelout<=1'b0;
18372: pixelout<=1'b0;
18373: pixelout<=1'b1;
18374: pixelout<=1'b1;
18375: pixelout<=1'b0;
18376: pixelout<=1'b1;
18377: pixelout<=1'b0;
18378: pixelout<=1'b1;
18379: pixelout<=1'b1;
18380: pixelout<=1'b0;
18381: pixelout<=1'b0;
18382: pixelout<=1'b0;
18383: pixelout<=1'b0;
18384: pixelout<=1'b0;
18385: pixelout<=1'b1;
18386: pixelout<=1'b1;
18387: pixelout<=1'b1;
18388: pixelout<=1'b1;
18389: pixelout<=1'b1;
18390: pixelout<=1'b1;
18391: pixelout<=1'b1;
18392: pixelout<=1'b1;
18393: pixelout<=1'b1;
18394: pixelout<=1'b1;
18395: pixelout<=1'b1;
18396: pixelout<=1'b0;
18397: pixelout<=1'b1;
18398: pixelout<=1'b0;
18399: pixelout<=1'b1;
18400: pixelout<=1'b1;
18401: pixelout<=1'b1;
18402: pixelout<=1'b0;
18403: pixelout<=1'b1;
18404: pixelout<=1'b0;
18405: pixelout<=1'b1;
18406: pixelout<=1'b1;
18407: pixelout<=1'b0;
18408: pixelout<=1'b1;
18409: pixelout<=1'b0;
18410: pixelout<=1'b0;
18411: pixelout<=1'b0;
18412: pixelout<=1'b0;
18413: pixelout<=1'b0;
18414: pixelout<=1'b1;
18415: pixelout<=1'b1;
18416: pixelout<=1'b1;
18417: pixelout<=1'b1;
18418: pixelout<=1'b0;
18419: pixelout<=1'b1;
18420: pixelout<=1'b0;
18421: pixelout<=1'b1;
18422: pixelout<=1'b0;
18423: pixelout<=1'b1;
18424: pixelout<=1'b0;
18425: pixelout<=1'b1;
18426: pixelout<=1'b1;
18427: pixelout<=1'b1;
18428: pixelout<=1'b0;
18429: pixelout<=1'b1;
18430: pixelout<=1'b0;
18431: pixelout<=1'b1;
18432: pixelout<=1'b1;
18433: pixelout<=1'b1;
18434: pixelout<=1'b1;
18435: pixelout<=1'b1;
18436: pixelout<=1'b1;
18437: pixelout<=1'b1;
18438: pixelout<=1'b1;
18439: pixelout<=1'b1;
18440: pixelout<=1'b1;
18441: pixelout<=1'b1;
18442: pixelout<=1'b1;
18443: pixelout<=1'b0;
18444: pixelout<=1'b1;
18445: pixelout<=1'b0;
18446: pixelout<=1'b0;
18447: pixelout<=1'b0;
18448: pixelout<=1'b0;
18449: pixelout<=1'b0;
18450: pixelout<=1'b1;
18451: pixelout<=1'b1;
18452: pixelout<=1'b0;
18453: pixelout<=1'b1;
18454: pixelout<=1'b0;
18455: pixelout<=1'b1;
18456: pixelout<=1'b1;
18457: pixelout<=1'b1;
18458: pixelout<=1'b0;
18459: pixelout<=1'b1;
18460: pixelout<=1'b0;
18461: pixelout<=1'b0;
18462: pixelout<=1'b0;
18463: pixelout<=1'b0;
18464: pixelout<=1'b0;
18465: pixelout<=1'b1;
18466: pixelout<=1'b1;
18467: pixelout<=1'b1;
18468: pixelout<=1'b1;
18469: pixelout<=1'b1;
18470: pixelout<=1'b1;
18471: pixelout<=1'b0;
18472: pixelout<=1'b1;
18473: pixelout<=1'b1;
18474: pixelout<=1'b1;
18475: pixelout<=1'b1;
18476: pixelout<=1'b1;
18477: pixelout<=1'b1;
18478: pixelout<=1'b1;
18479: pixelout<=1'b1;
18480: pixelout<=1'b1;
18481: pixelout<=1'b1;
18482: pixelout<=1'b1;
18483: pixelout<=1'b1;
18484: pixelout<=1'b1;
18485: pixelout<=1'b1;
18486: pixelout<=1'b1;
18487: pixelout<=1'b1;
18488: pixelout<=1'b1;
18489: pixelout<=1'b0;
18490: pixelout<=1'b1;
18491: pixelout<=1'b1;
18492: pixelout<=1'b1;
18493: pixelout<=1'b0;
18494: pixelout<=1'b1;
18495: pixelout<=1'b0;
18496: pixelout<=1'b1;
18497: pixelout<=1'b1;
18498: pixelout<=1'b1;
18499: pixelout<=1'b1;
18500: pixelout<=1'b1;
18501: pixelout<=1'b1;
18502: pixelout<=1'b1;
18503: pixelout<=1'b1;
18504: pixelout<=1'b1;
18505: pixelout<=1'b1;
18506: pixelout<=1'b1;
18507: pixelout<=1'b1;
18508: pixelout<=1'b0;
18509: pixelout<=1'b1;
18510: pixelout<=1'b0;
18511: pixelout<=1'b1;
18512: pixelout<=1'b1;
18513: pixelout<=1'b0;
18514: pixelout<=1'b1;
18515: pixelout<=1'b0;
18516: pixelout<=1'b1;
18517: pixelout<=1'b1;
18518: pixelout<=1'b0;
18519: pixelout<=1'b1;
18520: pixelout<=1'b1;
18521: pixelout<=1'b1;
18522: pixelout<=1'b1;
18523: pixelout<=1'b1;
18524: pixelout<=1'b0;
18525: pixelout<=1'b1;
18526: pixelout<=1'b1;
18527: pixelout<=1'b1;
18528: pixelout<=1'b1;
18529: pixelout<=1'b1;
18530: pixelout<=1'b1;
18531: pixelout<=1'b0;
18532: pixelout<=1'b1;
18533: pixelout<=1'b0;
18534: pixelout<=1'b1;
18535: pixelout<=1'b1;
18536: pixelout<=1'b1;
18537: pixelout<=1'b0;
18538: pixelout<=1'b1;
18539: pixelout<=1'b0;
18540: pixelout<=1'b1;
18541: pixelout<=1'b1;
18542: pixelout<=1'b0;
18543: pixelout<=1'b0;
18544: pixelout<=1'b1;
18545: pixelout<=1'b0;
18546: pixelout<=1'b0;
18547: pixelout<=1'b1;
18548: pixelout<=1'b1;
18549: pixelout<=1'b1;
18550: pixelout<=1'b0;
18551: pixelout<=1'b1;
18552: pixelout<=1'b1;
18553: pixelout<=1'b1;
18554: pixelout<=1'b1;
18555: pixelout<=1'b1;
18556: pixelout<=1'b1;
18557: pixelout<=1'b1;
18558: pixelout<=1'b1;
18559: pixelout<=1'b1;
18560: pixelout<=1'b1;
18561: pixelout<=1'b0;
18562: pixelout<=1'b1;
18563: pixelout<=1'b1;
18564: pixelout<=1'b1;
18565: pixelout<=1'b1;
18566: pixelout<=1'b1;
18567: pixelout<=1'b0;
18568: pixelout<=1'b1;
18569: pixelout<=1'b1;
18570: pixelout<=1'b1;
18571: pixelout<=1'b0;
18572: pixelout<=1'b1;
18573: pixelout<=1'b1;
18574: pixelout<=1'b0;
18575: pixelout<=1'b0;
18576: pixelout<=1'b1;
18577: pixelout<=1'b1;
18578: pixelout<=1'b1;
18579: pixelout<=1'b1;
18580: pixelout<=1'b1;
18581: pixelout<=1'b0;
18582: pixelout<=1'b1;
18583: pixelout<=1'b0;
18584: pixelout<=1'b0;
18585: pixelout<=1'b1;
18586: pixelout<=1'b1;
18587: pixelout<=1'b1;
18588: pixelout<=1'b0;
18589: pixelout<=1'b1;
18590: pixelout<=1'b1;
18591: pixelout<=1'b0;
18592: pixelout<=1'b0;
18593: pixelout<=1'b1;
18594: pixelout<=1'b0;
18595: pixelout<=1'b1;
18596: pixelout<=1'b1;
18597: pixelout<=1'b0;
18598: pixelout<=1'b1;
18599: pixelout<=1'b0;
18600: pixelout<=1'b1;
18601: pixelout<=1'b1;
18602: pixelout<=1'b1;
18603: pixelout<=1'b1;
18604: pixelout<=1'b1;
18605: pixelout<=1'b1;
18606: pixelout<=1'b1;
18607: pixelout<=1'b1;
18608: pixelout<=1'b0;
18609: pixelout<=1'b1;
18610: pixelout<=1'b1;
18611: pixelout<=1'b1;
18612: pixelout<=1'b1;
18613: pixelout<=1'b1;
18614: pixelout<=1'b1;
18615: pixelout<=1'b0;
18616: pixelout<=1'b1;
18617: pixelout<=1'b0;
18618: pixelout<=1'b1;
18619: pixelout<=1'b1;
18620: pixelout<=1'b0;
18621: pixelout<=1'b1;
18622: pixelout<=1'b1;
18623: pixelout<=1'b1;
18624: pixelout<=1'b1;
18625: pixelout<=1'b1;
18626: pixelout<=1'b1;
18627: pixelout<=1'b1;
18628: pixelout<=1'b1;
18629: pixelout<=1'b1;
18630: pixelout<=1'b1;
18631: pixelout<=1'b1;
18632: pixelout<=1'b1;
18633: pixelout<=1'b1;
18634: pixelout<=1'b1;
18635: pixelout<=1'b1;
18636: pixelout<=1'b0;
18637: pixelout<=1'b1;
18638: pixelout<=1'b0;
18639: pixelout<=1'b1;
18640: pixelout<=1'b1;
18641: pixelout<=1'b1;
18642: pixelout<=1'b0;
18643: pixelout<=1'b1;
18644: pixelout<=1'b0;
18645: pixelout<=1'b1;
18646: pixelout<=1'b1;
18647: pixelout<=1'b0;
18648: pixelout<=1'b1;
18649: pixelout<=1'b0;
18650: pixelout<=1'b1;
18651: pixelout<=1'b1;
18652: pixelout<=1'b1;
18653: pixelout<=1'b1;
18654: pixelout<=1'b1;
18655: pixelout<=1'b1;
18656: pixelout<=1'b1;
18657: pixelout<=1'b1;
18658: pixelout<=1'b0;
18659: pixelout<=1'b1;
18660: pixelout<=1'b0;
18661: pixelout<=1'b1;
18662: pixelout<=1'b0;
18663: pixelout<=1'b1;
18664: pixelout<=1'b0;
18665: pixelout<=1'b1;
18666: pixelout<=1'b1;
18667: pixelout<=1'b1;
18668: pixelout<=1'b0;
18669: pixelout<=1'b1;
18670: pixelout<=1'b0;
18671: pixelout<=1'b1;
18672: pixelout<=1'b1;
18673: pixelout<=1'b1;
18674: pixelout<=1'b1;
18675: pixelout<=1'b1;
18676: pixelout<=1'b1;
18677: pixelout<=1'b1;
18678: pixelout<=1'b1;
18679: pixelout<=1'b1;
18680: pixelout<=1'b1;
18681: pixelout<=1'b1;
18682: pixelout<=1'b1;
18683: pixelout<=1'b0;
18684: pixelout<=1'b1;
18685: pixelout<=1'b0;
18686: pixelout<=1'b1;
18687: pixelout<=1'b1;
18688: pixelout<=1'b1;
18689: pixelout<=1'b1;
18690: pixelout<=1'b1;
18691: pixelout<=1'b1;
18692: pixelout<=1'b0;
18693: pixelout<=1'b1;
18694: pixelout<=1'b0;
18695: pixelout<=1'b1;
18696: pixelout<=1'b1;
18697: pixelout<=1'b1;
18698: pixelout<=1'b0;
18699: pixelout<=1'b1;
18700: pixelout<=1'b0;
18701: pixelout<=1'b1;
18702: pixelout<=1'b1;
18703: pixelout<=1'b1;
18704: pixelout<=1'b1;
18705: pixelout<=1'b1;
18706: pixelout<=1'b1;
18707: pixelout<=1'b1;
18708: pixelout<=1'b1;
18709: pixelout<=1'b1;
18710: pixelout<=1'b1;
18711: pixelout<=1'b0;
18712: pixelout<=1'b1;
18713: pixelout<=1'b1;
18714: pixelout<=1'b1;
18715: pixelout<=1'b1;
18716: pixelout<=1'b1;
18717: pixelout<=1'b1;
18718: pixelout<=1'b1;
18719: pixelout<=1'b1;
18720: pixelout<=1'b1;
18721: pixelout<=1'b1;
18722: pixelout<=1'b1;
18723: pixelout<=1'b1;
18724: pixelout<=1'b1;
18725: pixelout<=1'b1;
18726: pixelout<=1'b1;
18727: pixelout<=1'b1;
18728: pixelout<=1'b1;
18729: pixelout<=1'b1;
18730: pixelout<=1'b0;
18731: pixelout<=1'b0;
18732: pixelout<=1'b0;
18733: pixelout<=1'b1;
18734: pixelout<=1'b1;
18735: pixelout<=1'b0;
18736: pixelout<=1'b1;
18737: pixelout<=1'b1;
18738: pixelout<=1'b1;
18739: pixelout<=1'b1;
18740: pixelout<=1'b1;
18741: pixelout<=1'b1;
18742: pixelout<=1'b1;
18743: pixelout<=1'b1;
18744: pixelout<=1'b1;
18745: pixelout<=1'b1;
18746: pixelout<=1'b1;
18747: pixelout<=1'b1;
18748: pixelout<=1'b0;
18749: pixelout<=1'b1;
18750: pixelout<=1'b0;
18751: pixelout<=1'b1;
18752: pixelout<=1'b1;
18753: pixelout<=1'b0;
18754: pixelout<=1'b1;
18755: pixelout<=1'b1;
18756: pixelout<=1'b0;
18757: pixelout<=1'b0;
18758: pixelout<=1'b1;
18759: pixelout<=1'b0;
18760: pixelout<=1'b1;
18761: pixelout<=1'b0;
18762: pixelout<=1'b0;
18763: pixelout<=1'b0;
18764: pixelout<=1'b0;
18765: pixelout<=1'b1;
18766: pixelout<=1'b1;
18767: pixelout<=1'b1;
18768: pixelout<=1'b1;
18769: pixelout<=1'b1;
18770: pixelout<=1'b1;
18771: pixelout<=1'b0;
18772: pixelout<=1'b1;
18773: pixelout<=1'b1;
18774: pixelout<=1'b0;
18775: pixelout<=1'b0;
18776: pixelout<=1'b0;
18777: pixelout<=1'b0;
18778: pixelout<=1'b1;
18779: pixelout<=1'b1;
18780: pixelout<=1'b0;
18781: pixelout<=1'b0;
18782: pixelout<=1'b1;
18783: pixelout<=1'b0;
18784: pixelout<=1'b1;
18785: pixelout<=1'b0;
18786: pixelout<=1'b0;
18787: pixelout<=1'b1;
18788: pixelout<=1'b1;
18789: pixelout<=1'b1;
18790: pixelout<=1'b1;
18791: pixelout<=1'b0;
18792: pixelout<=1'b0;
18793: pixelout<=1'b0;
18794: pixelout<=1'b1;
18795: pixelout<=1'b1;
18796: pixelout<=1'b1;
18797: pixelout<=1'b1;
18798: pixelout<=1'b1;
18799: pixelout<=1'b1;
18800: pixelout<=1'b1;
18801: pixelout<=1'b0;
18802: pixelout<=1'b1;
18803: pixelout<=1'b1;
18804: pixelout<=1'b1;
18805: pixelout<=1'b0;
18806: pixelout<=1'b0;
18807: pixelout<=1'b0;
18808: pixelout<=1'b0;
18809: pixelout<=1'b0;
18810: pixelout<=1'b1;
18811: pixelout<=1'b1;
18812: pixelout<=1'b0;
18813: pixelout<=1'b0;
18814: pixelout<=1'b1;
18815: pixelout<=1'b1;
18816: pixelout<=1'b1;
18817: pixelout<=1'b1;
18818: pixelout<=1'b1;
18819: pixelout<=1'b1;
18820: pixelout<=1'b1;
18821: pixelout<=1'b0;
18822: pixelout<=1'b1;
18823: pixelout<=1'b0;
18824: pixelout<=1'b0;
18825: pixelout<=1'b1;
18826: pixelout<=1'b1;
18827: pixelout<=1'b1;
18828: pixelout<=1'b1;
18829: pixelout<=1'b0;
18830: pixelout<=1'b0;
18831: pixelout<=1'b1;
18832: pixelout<=1'b0;
18833: pixelout<=1'b1;
18834: pixelout<=1'b0;
18835: pixelout<=1'b1;
18836: pixelout<=1'b1;
18837: pixelout<=1'b0;
18838: pixelout<=1'b1;
18839: pixelout<=1'b1;
18840: pixelout<=1'b0;
18841: pixelout<=1'b0;
18842: pixelout<=1'b0;
18843: pixelout<=1'b0;
18844: pixelout<=1'b1;
18845: pixelout<=1'b1;
18846: pixelout<=1'b1;
18847: pixelout<=1'b1;
18848: pixelout<=1'b1;
18849: pixelout<=1'b0;
18850: pixelout<=1'b0;
18851: pixelout<=1'b0;
18852: pixelout<=1'b0;
18853: pixelout<=1'b1;
18854: pixelout<=1'b1;
18855: pixelout<=1'b1;
18856: pixelout<=1'b0;
18857: pixelout<=1'b1;
18858: pixelout<=1'b1;
18859: pixelout<=1'b1;
18860: pixelout<=1'b1;
18861: pixelout<=1'b0;
18862: pixelout<=1'b0;
18863: pixelout<=1'b0;
18864: pixelout<=1'b0;
18865: pixelout<=1'b1;
18866: pixelout<=1'b1;
18867: pixelout<=1'b1;
18868: pixelout<=1'b1;
18869: pixelout<=1'b1;
18870: pixelout<=1'b1;
18871: pixelout<=1'b1;
18872: pixelout<=1'b1;
18873: pixelout<=1'b0;
18874: pixelout<=1'b0;
18875: pixelout<=1'b0;
18876: pixelout<=1'b0;
18877: pixelout<=1'b1;
18878: pixelout<=1'b1;
18879: pixelout<=1'b0;
18880: pixelout<=1'b0;
18881: pixelout<=1'b0;
18882: pixelout<=1'b1;
18883: pixelout<=1'b1;
18884: pixelout<=1'b0;
18885: pixelout<=1'b1;
18886: pixelout<=1'b1;
18887: pixelout<=1'b0;
18888: pixelout<=1'b1;
18889: pixelout<=1'b1;
18890: pixelout<=1'b0;
18891: pixelout<=1'b0;
18892: pixelout<=1'b0;
18893: pixelout<=1'b0;
18894: pixelout<=1'b1;
18895: pixelout<=1'b1;
18896: pixelout<=1'b1;
18897: pixelout<=1'b1;
18898: pixelout<=1'b1;
18899: pixelout<=1'b0;
18900: pixelout<=1'b1;
18901: pixelout<=1'b0;
18902: pixelout<=1'b1;
18903: pixelout<=1'b1;
18904: pixelout<=1'b0;
18905: pixelout<=1'b1;
18906: pixelout<=1'b1;
18907: pixelout<=1'b1;
18908: pixelout<=1'b0;
18909: pixelout<=1'b1;
18910: pixelout<=1'b1;
18911: pixelout<=1'b0;
18912: pixelout<=1'b0;
18913: pixelout<=1'b0;
18914: pixelout<=1'b1;
18915: pixelout<=1'b1;
18916: pixelout<=1'b1;
18917: pixelout<=1'b1;
18918: pixelout<=1'b1;
18919: pixelout<=1'b1;
18920: pixelout<=1'b1;
18921: pixelout<=1'b1;
18922: pixelout<=1'b1;
18923: pixelout<=1'b0;
18924: pixelout<=1'b1;
18925: pixelout<=1'b1;
18926: pixelout<=1'b0;
18927: pixelout<=1'b0;
18928: pixelout<=1'b0;
18929: pixelout<=1'b0;
18930: pixelout<=1'b1;
18931: pixelout<=1'b1;
18932: pixelout<=1'b0;
18933: pixelout<=1'b1;
18934: pixelout<=1'b0;
18935: pixelout<=1'b0;
18936: pixelout<=1'b0;
18937: pixelout<=1'b0;
18938: pixelout<=1'b1;
18939: pixelout<=1'b1;
18940: pixelout<=1'b1;
18941: pixelout<=1'b0;
18942: pixelout<=1'b0;
18943: pixelout<=1'b0;
18944: pixelout<=1'b0;
18945: pixelout<=1'b1;
18946: pixelout<=1'b1;
18947: pixelout<=1'b1;
18948: pixelout<=1'b0;
18949: pixelout<=1'b0;
18950: pixelout<=1'b0;
18951: pixelout<=1'b0;
18952: pixelout<=1'b1;
18953: pixelout<=1'b1;
18954: pixelout<=1'b1;
18955: pixelout<=1'b1;
18956: pixelout<=1'b1;
18957: pixelout<=1'b1;
18958: pixelout<=1'b1;
18959: pixelout<=1'b1;
18960: pixelout<=1'b1;
18961: pixelout<=1'b1;
18962: pixelout<=1'b1;
18963: pixelout<=1'b1;
18964: pixelout<=1'b1;
18965: pixelout<=1'b1;
18966: pixelout<=1'b1;
18967: pixelout<=1'b1;
18968: pixelout<=1'b1;
18969: pixelout<=1'b1;
18970: pixelout<=1'b1;
18971: pixelout<=1'b1;
18972: pixelout<=1'b1;
18973: pixelout<=1'b1;
18974: pixelout<=1'b1;
18975: pixelout<=1'b1;
18976: pixelout<=1'b1;
18977: pixelout<=1'b1;
18978: pixelout<=1'b1;
18979: pixelout<=1'b1;
18980: pixelout<=1'b1;
18981: pixelout<=1'b1;
18982: pixelout<=1'b1;
18983: pixelout<=1'b1;
18984: pixelout<=1'b1;
18985: pixelout<=1'b1;
18986: pixelout<=1'b1;
18987: pixelout<=1'b1;
18988: pixelout<=1'b1;
18989: pixelout<=1'b1;
18990: pixelout<=1'b1;
18991: pixelout<=1'b1;
18992: pixelout<=1'b1;
18993: pixelout<=1'b1;
18994: pixelout<=1'b1;
18995: pixelout<=1'b1;
18996: pixelout<=1'b1;
18997: pixelout<=1'b1;
18998: pixelout<=1'b1;
18999: pixelout<=1'b1;
19000: pixelout<=1'b1;
19001: pixelout<=1'b1;
19002: pixelout<=1'b1;
19003: pixelout<=1'b1;
19004: pixelout<=1'b1;
19005: pixelout<=1'b1;
19006: pixelout<=1'b1;
19007: pixelout<=1'b1;
19008: pixelout<=1'b1;
19009: pixelout<=1'b1;
19010: pixelout<=1'b1;
19011: pixelout<=1'b1;
19012: pixelout<=1'b1;
19013: pixelout<=1'b1;
19014: pixelout<=1'b1;
19015: pixelout<=1'b1;
19016: pixelout<=1'b1;
19017: pixelout<=1'b0;
19018: pixelout<=1'b1;
19019: pixelout<=1'b1;
19020: pixelout<=1'b1;
19021: pixelout<=1'b1;
19022: pixelout<=1'b1;
19023: pixelout<=1'b1;
19024: pixelout<=1'b1;
19025: pixelout<=1'b1;
19026: pixelout<=1'b0;
19027: pixelout<=1'b1;
19028: pixelout<=1'b1;
19029: pixelout<=1'b1;
19030: pixelout<=1'b1;
19031: pixelout<=1'b1;
19032: pixelout<=1'b1;
19033: pixelout<=1'b1;
19034: pixelout<=1'b1;
19035: pixelout<=1'b1;
19036: pixelout<=1'b1;
19037: pixelout<=1'b1;
19038: pixelout<=1'b1;
19039: pixelout<=1'b1;
19040: pixelout<=1'b1;
19041: pixelout<=1'b1;
19042: pixelout<=1'b1;
19043: pixelout<=1'b1;
19044: pixelout<=1'b1;
19045: pixelout<=1'b1;
19046: pixelout<=1'b1;
19047: pixelout<=1'b1;
19048: pixelout<=1'b1;
19049: pixelout<=1'b1;
19050: pixelout<=1'b1;
19051: pixelout<=1'b1;
19052: pixelout<=1'b1;
19053: pixelout<=1'b1;
19054: pixelout<=1'b1;
19055: pixelout<=1'b1;
19056: pixelout<=1'b1;
19057: pixelout<=1'b1;
19058: pixelout<=1'b1;
19059: pixelout<=1'b1;
19060: pixelout<=1'b1;
19061: pixelout<=1'b1;
19062: pixelout<=1'b1;
19063: pixelout<=1'b1;
19064: pixelout<=1'b0;
19065: pixelout<=1'b1;
19066: pixelout<=1'b1;
19067: pixelout<=1'b1;
19068: pixelout<=1'b1;
19069: pixelout<=1'b1;
19070: pixelout<=1'b1;
19071: pixelout<=1'b1;
19072: pixelout<=1'b1;
19073: pixelout<=1'b1;
19074: pixelout<=1'b1;
19075: pixelout<=1'b1;
19076: pixelout<=1'b1;
19077: pixelout<=1'b1;
19078: pixelout<=1'b1;
19079: pixelout<=1'b1;
19080: pixelout<=1'b1;
19081: pixelout<=1'b1;
19082: pixelout<=1'b1;
19083: pixelout<=1'b1;
19084: pixelout<=1'b1;
19085: pixelout<=1'b1;
19086: pixelout<=1'b1;
19087: pixelout<=1'b1;
19088: pixelout<=1'b1;
19089: pixelout<=1'b1;
19090: pixelout<=1'b1;
19091: pixelout<=1'b1;
19092: pixelout<=1'b1;
19093: pixelout<=1'b1;
19094: pixelout<=1'b1;
19095: pixelout<=1'b1;
19096: pixelout<=1'b1;
19097: pixelout<=1'b1;
19098: pixelout<=1'b1;
19099: pixelout<=1'b1;
19100: pixelout<=1'b1;
19101: pixelout<=1'b1;
19102: pixelout<=1'b1;
19103: pixelout<=1'b1;
19104: pixelout<=1'b1;
19105: pixelout<=1'b1;
19106: pixelout<=1'b1;
19107: pixelout<=1'b1;
19108: pixelout<=1'b1;
19109: pixelout<=1'b1;
19110: pixelout<=1'b1;
19111: pixelout<=1'b1;
19112: pixelout<=1'b1;
19113: pixelout<=1'b1;
19114: pixelout<=1'b1;
19115: pixelout<=1'b1;
19116: pixelout<=1'b0;
19117: pixelout<=1'b1;
19118: pixelout<=1'b1;
19119: pixelout<=1'b1;
19120: pixelout<=1'b1;
19121: pixelout<=1'b1;
19122: pixelout<=1'b1;
19123: pixelout<=1'b1;
19124: pixelout<=1'b1;
19125: pixelout<=1'b1;
19126: pixelout<=1'b1;
19127: pixelout<=1'b1;
19128: pixelout<=1'b1;
19129: pixelout<=1'b1;
19130: pixelout<=1'b1;
19131: pixelout<=1'b1;
19132: pixelout<=1'b1;
19133: pixelout<=1'b1;
19134: pixelout<=1'b1;
19135: pixelout<=1'b1;
19136: pixelout<=1'b1;
19137: pixelout<=1'b1;
19138: pixelout<=1'b1;
19139: pixelout<=1'b1;
19140: pixelout<=1'b1;
19141: pixelout<=1'b1;
19142: pixelout<=1'b1;
19143: pixelout<=1'b1;
19144: pixelout<=1'b1;
19145: pixelout<=1'b1;
19146: pixelout<=1'b1;
19147: pixelout<=1'b1;
19148: pixelout<=1'b1;
19149: pixelout<=1'b1;
19150: pixelout<=1'b1;
19151: pixelout<=1'b1;
19152: pixelout<=1'b1;
19153: pixelout<=1'b1;
19154: pixelout<=1'b1;
19155: pixelout<=1'b1;
19156: pixelout<=1'b1;
19157: pixelout<=1'b1;
19158: pixelout<=1'b1;
19159: pixelout<=1'b1;
19160: pixelout<=1'b1;
19161: pixelout<=1'b1;
19162: pixelout<=1'b1;
19163: pixelout<=1'b1;
19164: pixelout<=1'b1;
19165: pixelout<=1'b1;
19166: pixelout<=1'b1;
19167: pixelout<=1'b1;
19168: pixelout<=1'b1;
19169: pixelout<=1'b1;
19170: pixelout<=1'b1;
19171: pixelout<=1'b1;
19172: pixelout<=1'b1;
19173: pixelout<=1'b1;
19174: pixelout<=1'b0;
19175: pixelout<=1'b1;
19176: pixelout<=1'b1;
19177: pixelout<=1'b1;
19178: pixelout<=1'b1;
19179: pixelout<=1'b1;
19180: pixelout<=1'b1;
19181: pixelout<=1'b1;
19182: pixelout<=1'b1;
19183: pixelout<=1'b1;
19184: pixelout<=1'b1;
19185: pixelout<=1'b1;
19186: pixelout<=1'b1;
19187: pixelout<=1'b1;
19188: pixelout<=1'b1;
19189: pixelout<=1'b1;
19190: pixelout<=1'b1;
19191: pixelout<=1'b1;
19192: pixelout<=1'b1;
19193: pixelout<=1'b1;
19194: pixelout<=1'b1;
19195: pixelout<=1'b1;
19196: pixelout<=1'b1;
19197: pixelout<=1'b1;
19198: pixelout<=1'b1;
19199: pixelout<=1'b1;
19200: pixelout<=1'b1;
19201: pixelout<=1'b1;
19202: pixelout<=1'b1;
19203: pixelout<=1'b1;
19204: pixelout<=1'b1;
19205: pixelout<=1'b1;
19206: pixelout<=1'b1;
19207: pixelout<=1'b1;
19208: pixelout<=1'b1;
19209: pixelout<=1'b1;
19210: pixelout<=1'b1;
19211: pixelout<=1'b1;
19212: pixelout<=1'b1;
19213: pixelout<=1'b1;
19214: pixelout<=1'b1;
19215: pixelout<=1'b1;
19216: pixelout<=1'b1;
19217: pixelout<=1'b1;
19218: pixelout<=1'b1;
19219: pixelout<=1'b1;
19220: pixelout<=1'b1;
19221: pixelout<=1'b1;
19222: pixelout<=1'b1;
19223: pixelout<=1'b1;
19224: pixelout<=1'b1;
19225: pixelout<=1'b1;
19226: pixelout<=1'b1;
19227: pixelout<=1'b1;
19228: pixelout<=1'b1;
19229: pixelout<=1'b1;
19230: pixelout<=1'b1;
19231: pixelout<=1'b1;
19232: pixelout<=1'b1;
19233: pixelout<=1'b1;
19234: pixelout<=1'b1;
19235: pixelout<=1'b1;
19236: pixelout<=1'b1;
19237: pixelout<=1'b1;
19238: pixelout<=1'b1;
19239: pixelout<=1'b1;
19240: pixelout<=1'b1;
19241: pixelout<=1'b1;
19242: pixelout<=1'b1;
19243: pixelout<=1'b1;
19244: pixelout<=1'b1;
19245: pixelout<=1'b1;
19246: pixelout<=1'b1;
19247: pixelout<=1'b1;
19248: pixelout<=1'b1;
19249: pixelout<=1'b1;
19250: pixelout<=1'b1;
19251: pixelout<=1'b1;
19252: pixelout<=1'b1;
19253: pixelout<=1'b0;
19254: pixelout<=1'b0;
19255: pixelout<=1'b0;
19256: pixelout<=1'b0;
19257: pixelout<=1'b1;
19258: pixelout<=1'b1;
19259: pixelout<=1'b1;
19260: pixelout<=1'b1;
19261: pixelout<=1'b1;
19262: pixelout<=1'b1;
19263: pixelout<=1'b1;
19264: pixelout<=1'b1;
19265: pixelout<=1'b0;
19266: pixelout<=1'b1;
19267: pixelout<=1'b1;
19268: pixelout<=1'b1;
19269: pixelout<=1'b1;
19270: pixelout<=1'b1;
19271: pixelout<=1'b1;
19272: pixelout<=1'b1;
19273: pixelout<=1'b1;
19274: pixelout<=1'b1;
19275: pixelout<=1'b1;
19276: pixelout<=1'b1;
19277: pixelout<=1'b1;
19278: pixelout<=1'b1;
19279: pixelout<=1'b1;
19280: pixelout<=1'b1;
19281: pixelout<=1'b1;
19282: pixelout<=1'b1;
19283: pixelout<=1'b1;
19284: pixelout<=1'b1;
19285: pixelout<=1'b1;
19286: pixelout<=1'b1;
19287: pixelout<=1'b1;
19288: pixelout<=1'b1;
19289: pixelout<=1'b1;
19290: pixelout<=1'b1;
19291: pixelout<=1'b1;
19292: pixelout<=1'b1;
19293: pixelout<=1'b1;
19294: pixelout<=1'b1;
19295: pixelout<=1'b1;
19296: pixelout<=1'b1;
19297: pixelout<=1'b1;
19298: pixelout<=1'b1;
19299: pixelout<=1'b1;
19300: pixelout<=1'b1;
19301: pixelout<=1'b1;
19302: pixelout<=1'b1;
19303: pixelout<=1'b0;
19304: pixelout<=1'b1;
19305: pixelout<=1'b1;
19306: pixelout<=1'b1;
19307: pixelout<=1'b1;
19308: pixelout<=1'b1;
19309: pixelout<=1'b1;
19310: pixelout<=1'b1;
19311: pixelout<=1'b1;
19312: pixelout<=1'b1;
19313: pixelout<=1'b1;
19314: pixelout<=1'b1;
19315: pixelout<=1'b1;
19316: pixelout<=1'b1;
19317: pixelout<=1'b1;
19318: pixelout<=1'b1;
19319: pixelout<=1'b1;
19320: pixelout<=1'b1;
19321: pixelout<=1'b1;
19322: pixelout<=1'b1;
19323: pixelout<=1'b1;
19324: pixelout<=1'b1;
19325: pixelout<=1'b1;
19326: pixelout<=1'b1;
19327: pixelout<=1'b1;
19328: pixelout<=1'b1;
19329: pixelout<=1'b1;
19330: pixelout<=1'b1;
19331: pixelout<=1'b1;
19332: pixelout<=1'b1;
19333: pixelout<=1'b1;
19334: pixelout<=1'b1;
19335: pixelout<=1'b1;
19336: pixelout<=1'b1;
19337: pixelout<=1'b1;
19338: pixelout<=1'b1;
19339: pixelout<=1'b1;
19340: pixelout<=1'b1;
19341: pixelout<=1'b1;
19342: pixelout<=1'b1;
19343: pixelout<=1'b1;
19344: pixelout<=1'b1;
19345: pixelout<=1'b1;
19346: pixelout<=1'b1;
19347: pixelout<=1'b1;
19348: pixelout<=1'b1;
19349: pixelout<=1'b1;
19350: pixelout<=1'b1;
19351: pixelout<=1'b1;
19352: pixelout<=1'b0;
19353: pixelout<=1'b0;
19354: pixelout<=1'b0;
19355: pixelout<=1'b0;
19356: pixelout<=1'b1;
19357: pixelout<=1'b1;
19358: pixelout<=1'b1;
19359: pixelout<=1'b1;
19360: pixelout<=1'b1;
19361: pixelout<=1'b1;
19362: pixelout<=1'b1;
19363: pixelout<=1'b1;
19364: pixelout<=1'b1;
19365: pixelout<=1'b1;
19366: pixelout<=1'b1;
19367: pixelout<=1'b1;
19368: pixelout<=1'b1;
19369: pixelout<=1'b1;
19370: pixelout<=1'b1;
19371: pixelout<=1'b1;
19372: pixelout<=1'b1;
19373: pixelout<=1'b1;
19374: pixelout<=1'b1;
19375: pixelout<=1'b1;
19376: pixelout<=1'b1;
19377: pixelout<=1'b1;
19378: pixelout<=1'b1;
19379: pixelout<=1'b1;
19380: pixelout<=1'b1;
19381: pixelout<=1'b1;
19382: pixelout<=1'b1;
19383: pixelout<=1'b1;
19384: pixelout<=1'b1;
19385: pixelout<=1'b1;
19386: pixelout<=1'b1;
19387: pixelout<=1'b1;
19388: pixelout<=1'b1;
19389: pixelout<=1'b1;
19390: pixelout<=1'b1;
19391: pixelout<=1'b1;
19392: pixelout<=1'b1;
19393: pixelout<=1'b1;
19394: pixelout<=1'b1;
19395: pixelout<=1'b1;
19396: pixelout<=1'b1;
19397: pixelout<=1'b1;
19398: pixelout<=1'b1;
19399: pixelout<=1'b1;
19400: pixelout<=1'b1;
19401: pixelout<=1'b1;
19402: pixelout<=1'b1;
19403: pixelout<=1'b1;
19404: pixelout<=1'b1;
19405: pixelout<=1'b1;
19406: pixelout<=1'b1;
19407: pixelout<=1'b1;
19408: pixelout<=1'b1;
19409: pixelout<=1'b1;
19410: pixelout<=1'b1;
19411: pixelout<=1'b1;
19412: pixelout<=1'b1;
19413: pixelout<=1'b1;
19414: pixelout<=1'b0;
19415: pixelout<=1'b1;
19416: pixelout<=1'b1;
19417: pixelout<=1'b1;
19418: pixelout<=1'b1;
19419: pixelout<=1'b1;
19420: pixelout<=1'b1;
19421: pixelout<=1'b1;
19422: pixelout<=1'b1;
19423: pixelout<=1'b1;
19424: pixelout<=1'b1;
19425: pixelout<=1'b1;
19426: pixelout<=1'b1;
19427: pixelout<=1'b1;
19428: pixelout<=1'b1;
19429: pixelout<=1'b1;
19430: pixelout<=1'b1;
19431: pixelout<=1'b1;
19432: pixelout<=1'b1;
19433: pixelout<=1'b1;
19434: pixelout<=1'b1;
19435: pixelout<=1'b1;
19436: pixelout<=1'b1;
19437: pixelout<=1'b1;
19438: pixelout<=1'b1;
19439: pixelout<=1'b1;
19440: pixelout<=1'b1;
19441: pixelout<=1'b1;
19442: pixelout<=1'b1;
19443: pixelout<=1'b1;
19444: pixelout<=1'b1;
19445: pixelout<=1'b1;
19446: pixelout<=1'b1;
19447: pixelout<=1'b1;
19448: pixelout<=1'b1;
19449: pixelout<=1'b1;
19450: pixelout<=1'b1;
19451: pixelout<=1'b1;
19452: pixelout<=1'b1;
19453: pixelout<=1'b1;
19454: pixelout<=1'b1;
19455: pixelout<=1'b1;
19456: pixelout<=1'b1;
19457: pixelout<=1'b1;
19458: pixelout<=1'b1;
19459: pixelout<=1'b1;
19460: pixelout<=1'b1;
19461: pixelout<=1'b1;
19462: pixelout<=1'b1;
19463: pixelout<=1'b1;
19464: pixelout<=1'b1;
19465: pixelout<=1'b1;
19466: pixelout<=1'b1;
19467: pixelout<=1'b1;
19468: pixelout<=1'b1;
19469: pixelout<=1'b1;
19470: pixelout<=1'b1;
19471: pixelout<=1'b1;
19472: pixelout<=1'b1;
19473: pixelout<=1'b1;
19474: pixelout<=1'b1;
19475: pixelout<=1'b1;
19476: pixelout<=1'b1;
19477: pixelout<=1'b1;
19478: pixelout<=1'b1;
19479: pixelout<=1'b1;
19480: pixelout<=1'b1;
19481: pixelout<=1'b1;
19482: pixelout<=1'b1;
19483: pixelout<=1'b1;
19484: pixelout<=1'b1;
19485: pixelout<=1'b1;
19486: pixelout<=1'b1;
19487: pixelout<=1'b1;
19488: pixelout<=1'b1;
19489: pixelout<=1'b1;
19490: pixelout<=1'b1;
19491: pixelout<=1'b1;
19492: pixelout<=1'b1;
19493: pixelout<=1'b1;
19494: pixelout<=1'b1;
19495: pixelout<=1'b1;
19496: pixelout<=1'b1;
19497: pixelout<=1'b1;
19498: pixelout<=1'b1;
19499: pixelout<=1'b1;
19500: pixelout<=1'b1;
19501: pixelout<=1'b1;
19502: pixelout<=1'b1;
19503: pixelout<=1'b1;
19504: pixelout<=1'b1;
19505: pixelout<=1'b1;
19506: pixelout<=1'b1;
19507: pixelout<=1'b1;
19508: pixelout<=1'b1;
19509: pixelout<=1'b1;
19510: pixelout<=1'b1;
19511: pixelout<=1'b1;
19512: pixelout<=1'b1;
19513: pixelout<=1'b1;
19514: pixelout<=1'b1;
19515: pixelout<=1'b1;
19516: pixelout<=1'b1;
19517: pixelout<=1'b1;
19518: pixelout<=1'b1;
19519: pixelout<=1'b1;
19520: pixelout<=1'b1;
19521: pixelout<=1'b1;
19522: pixelout<=1'b1;
19523: pixelout<=1'b1;
19524: pixelout<=1'b1;
19525: pixelout<=1'b1;
19526: pixelout<=1'b1;
19527: pixelout<=1'b1;
19528: pixelout<=1'b1;
19529: pixelout<=1'b1;
19530: pixelout<=1'b1;
19531: pixelout<=1'b1;
19532: pixelout<=1'b1;
19533: pixelout<=1'b1;
19534: pixelout<=1'b1;
19535: pixelout<=1'b1;
19536: pixelout<=1'b1;
19537: pixelout<=1'b1;
19538: pixelout<=1'b1;
19539: pixelout<=1'b1;
19540: pixelout<=1'b1;
19541: pixelout<=1'b1;
19542: pixelout<=1'b1;
19543: pixelout<=1'b1;
19544: pixelout<=1'b1;
19545: pixelout<=1'b1;
19546: pixelout<=1'b1;
19547: pixelout<=1'b1;
19548: pixelout<=1'b1;
19549: pixelout<=1'b1;
19550: pixelout<=1'b1;
19551: pixelout<=1'b1;
19552: pixelout<=1'b1;
19553: pixelout<=1'b1;
19554: pixelout<=1'b1;
19555: pixelout<=1'b1;
19556: pixelout<=1'b1;
19557: pixelout<=1'b1;
19558: pixelout<=1'b1;
19559: pixelout<=1'b1;
19560: pixelout<=1'b1;
19561: pixelout<=1'b1;
19562: pixelout<=1'b1;
19563: pixelout<=1'b1;
19564: pixelout<=1'b1;
19565: pixelout<=1'b1;
19566: pixelout<=1'b1;
19567: pixelout<=1'b1;
19568: pixelout<=1'b1;
19569: pixelout<=1'b1;
19570: pixelout<=1'b1;
19571: pixelout<=1'b1;
19572: pixelout<=1'b1;
19573: pixelout<=1'b1;
19574: pixelout<=1'b1;
19575: pixelout<=1'b1;
19576: pixelout<=1'b1;
19577: pixelout<=1'b1;
19578: pixelout<=1'b1;
19579: pixelout<=1'b1;
19580: pixelout<=1'b1;
19581: pixelout<=1'b1;
19582: pixelout<=1'b1;
19583: pixelout<=1'b1;
19584: pixelout<=1'b1;
19585: pixelout<=1'b1;
19586: pixelout<=1'b1;
19587: pixelout<=1'b1;
19588: pixelout<=1'b1;
19589: pixelout<=1'b1;
19590: pixelout<=1'b1;
19591: pixelout<=1'b1;
19592: pixelout<=1'b1;
19593: pixelout<=1'b1;
19594: pixelout<=1'b1;
19595: pixelout<=1'b1;
19596: pixelout<=1'b1;
19597: pixelout<=1'b1;
19598: pixelout<=1'b1;
19599: pixelout<=1'b1;
19600: pixelout<=1'b1;
19601: pixelout<=1'b1;
19602: pixelout<=1'b1;
19603: pixelout<=1'b1;
19604: pixelout<=1'b1;
19605: pixelout<=1'b1;
19606: pixelout<=1'b1;
19607: pixelout<=1'b1;
19608: pixelout<=1'b1;
19609: pixelout<=1'b1;
19610: pixelout<=1'b1;
19611: pixelout<=1'b1;
19612: pixelout<=1'b1;
19613: pixelout<=1'b1;
19614: pixelout<=1'b1;
19615: pixelout<=1'b1;
19616: pixelout<=1'b1;
19617: pixelout<=1'b1;
19618: pixelout<=1'b1;
19619: pixelout<=1'b1;
19620: pixelout<=1'b1;
19621: pixelout<=1'b1;
19622: pixelout<=1'b1;
19623: pixelout<=1'b1;
19624: pixelout<=1'b1;
19625: pixelout<=1'b1;
19626: pixelout<=1'b1;
19627: pixelout<=1'b1;
19628: pixelout<=1'b1;
19629: pixelout<=1'b1;
19630: pixelout<=1'b1;
19631: pixelout<=1'b1;
19632: pixelout<=1'b1;
19633: pixelout<=1'b1;
19634: pixelout<=1'b1;
19635: pixelout<=1'b1;
19636: pixelout<=1'b1;
19637: pixelout<=1'b1;
19638: pixelout<=1'b1;
19639: pixelout<=1'b1;
19640: pixelout<=1'b1;
19641: pixelout<=1'b1;
19642: pixelout<=1'b1;
19643: pixelout<=1'b1;
19644: pixelout<=1'b1;
19645: pixelout<=1'b1;
19646: pixelout<=1'b1;
19647: pixelout<=1'b1;
19648: pixelout<=1'b1;
19649: pixelout<=1'b1;
19650: pixelout<=1'b1;
19651: pixelout<=1'b1;
19652: pixelout<=1'b1;
19653: pixelout<=1'b1;
19654: pixelout<=1'b1;
19655: pixelout<=1'b1;
19656: pixelout<=1'b1;
19657: pixelout<=1'b1;
19658: pixelout<=1'b1;
19659: pixelout<=1'b1;
19660: pixelout<=1'b1;
19661: pixelout<=1'b1;
19662: pixelout<=1'b1;
19663: pixelout<=1'b1;
19664: pixelout<=1'b1;
19665: pixelout<=1'b1;
19666: pixelout<=1'b1;
19667: pixelout<=1'b1;
19668: pixelout<=1'b1;
19669: pixelout<=1'b1;
19670: pixelout<=1'b1;
19671: pixelout<=1'b1;
19672: pixelout<=1'b1;
19673: pixelout<=1'b1;
19674: pixelout<=1'b1;
19675: pixelout<=1'b1;
19676: pixelout<=1'b1;
19677: pixelout<=1'b1;
19678: pixelout<=1'b1;
19679: pixelout<=1'b1;
19680: pixelout<=1'b1;
19681: pixelout<=1'b1;
19682: pixelout<=1'b1;
19683: pixelout<=1'b1;
19684: pixelout<=1'b1;
19685: pixelout<=1'b1;
19686: pixelout<=1'b1;
19687: pixelout<=1'b1;
19688: pixelout<=1'b1;
19689: pixelout<=1'b1;
19690: pixelout<=1'b1;
19691: pixelout<=1'b1;
19692: pixelout<=1'b1;
19693: pixelout<=1'b1;
19694: pixelout<=1'b1;
19695: pixelout<=1'b1;
19696: pixelout<=1'b1;
19697: pixelout<=1'b1;
19698: pixelout<=1'b1;
19699: pixelout<=1'b1;
19700: pixelout<=1'b1;
19701: pixelout<=1'b1;
19702: pixelout<=1'b1;
19703: pixelout<=1'b1;
19704: pixelout<=1'b1;
19705: pixelout<=1'b1;
19706: pixelout<=1'b1;
19707: pixelout<=1'b1;
19708: pixelout<=1'b1;
19709: pixelout<=1'b1;
19710: pixelout<=1'b1;
19711: pixelout<=1'b1;
19712: pixelout<=1'b1;
19713: pixelout<=1'b1;
19714: pixelout<=1'b1;
19715: pixelout<=1'b1;
19716: pixelout<=1'b1;
19717: pixelout<=1'b1;
19718: pixelout<=1'b1;
19719: pixelout<=1'b1;
19720: pixelout<=1'b1;
19721: pixelout<=1'b1;
19722: pixelout<=1'b1;
19723: pixelout<=1'b1;
19724: pixelout<=1'b1;
19725: pixelout<=1'b1;
19726: pixelout<=1'b1;
19727: pixelout<=1'b1;
19728: pixelout<=1'b1;
19729: pixelout<=1'b1;
19730: pixelout<=1'b1;
19731: pixelout<=1'b1;
19732: pixelout<=1'b1;
19733: pixelout<=1'b1;
19734: pixelout<=1'b1;
19735: pixelout<=1'b1;
19736: pixelout<=1'b1;
19737: pixelout<=1'b1;
19738: pixelout<=1'b1;
19739: pixelout<=1'b1;
19740: pixelout<=1'b1;
19741: pixelout<=1'b1;
19742: pixelout<=1'b1;
19743: pixelout<=1'b1;
19744: pixelout<=1'b1;
19745: pixelout<=1'b1;
19746: pixelout<=1'b1;
19747: pixelout<=1'b1;
19748: pixelout<=1'b1;
19749: pixelout<=1'b1;
19750: pixelout<=1'b1;
19751: pixelout<=1'b1;
19752: pixelout<=1'b1;
19753: pixelout<=1'b1;
19754: pixelout<=1'b1;
19755: pixelout<=1'b1;
19756: pixelout<=1'b1;
19757: pixelout<=1'b1;
19758: pixelout<=1'b1;
19759: pixelout<=1'b1;
19760: pixelout<=1'b1;
19761: pixelout<=1'b1;
19762: pixelout<=1'b1;
19763: pixelout<=1'b1;
19764: pixelout<=1'b1;
19765: pixelout<=1'b1;
19766: pixelout<=1'b1;
19767: pixelout<=1'b1;
19768: pixelout<=1'b1;
19769: pixelout<=1'b1;
19770: pixelout<=1'b1;
19771: pixelout<=1'b1;
19772: pixelout<=1'b1;
19773: pixelout<=1'b1;
19774: pixelout<=1'b1;
19775: pixelout<=1'b1;
19776: pixelout<=1'b1;
19777: pixelout<=1'b1;
19778: pixelout<=1'b1;
19779: pixelout<=1'b1;
19780: pixelout<=1'b1;
19781: pixelout<=1'b1;
19782: pixelout<=1'b1;
19783: pixelout<=1'b1;
19784: pixelout<=1'b1;
19785: pixelout<=1'b1;
19786: pixelout<=1'b1;
19787: pixelout<=1'b1;
19788: pixelout<=1'b1;
19789: pixelout<=1'b1;
19790: pixelout<=1'b1;
19791: pixelout<=1'b1;
19792: pixelout<=1'b1;
19793: pixelout<=1'b1;
19794: pixelout<=1'b1;
19795: pixelout<=1'b1;
19796: pixelout<=1'b1;
19797: pixelout<=1'b1;
19798: pixelout<=1'b1;
19799: pixelout<=1'b1;
19800: pixelout<=1'b1;
19801: pixelout<=1'b1;
19802: pixelout<=1'b1;
19803: pixelout<=1'b1;
19804: pixelout<=1'b1;
19805: pixelout<=1'b1;
19806: pixelout<=1'b1;
19807: pixelout<=1'b1;
19808: pixelout<=1'b1;
19809: pixelout<=1'b1;
19810: pixelout<=1'b1;
19811: pixelout<=1'b1;
19812: pixelout<=1'b1;
19813: pixelout<=1'b1;
19814: pixelout<=1'b1;
19815: pixelout<=1'b1;
19816: pixelout<=1'b1;
19817: pixelout<=1'b1;
19818: pixelout<=1'b1;
19819: pixelout<=1'b1;
19820: pixelout<=1'b1;
19821: pixelout<=1'b1;
19822: pixelout<=1'b1;
19823: pixelout<=1'b1;
19824: pixelout<=1'b1;
19825: pixelout<=1'b1;
19826: pixelout<=1'b1;
19827: pixelout<=1'b1;
19828: pixelout<=1'b1;
19829: pixelout<=1'b1;
19830: pixelout<=1'b1;
19831: pixelout<=1'b1;
19832: pixelout<=1'b1;
19833: pixelout<=1'b1;
19834: pixelout<=1'b1;
19835: pixelout<=1'b1;
19836: pixelout<=1'b1;
19837: pixelout<=1'b1;
19838: pixelout<=1'b1;
19839: pixelout<=1'b1;
19840: pixelout<=1'b1;
19841: pixelout<=1'b1;
19842: pixelout<=1'b1;
19843: pixelout<=1'b1;
19844: pixelout<=1'b1;
19845: pixelout<=1'b1;
19846: pixelout<=1'b1;
19847: pixelout<=1'b1;
19848: pixelout<=1'b1;
19849: pixelout<=1'b1;
19850: pixelout<=1'b1;
19851: pixelout<=1'b1;
19852: pixelout<=1'b1;
19853: pixelout<=1'b1;
19854: pixelout<=1'b1;
19855: pixelout<=1'b1;
19856: pixelout<=1'b1;
19857: pixelout<=1'b1;
19858: pixelout<=1'b1;
19859: pixelout<=1'b1;
19860: pixelout<=1'b1;
19861: pixelout<=1'b1;
19862: pixelout<=1'b1;
19863: pixelout<=1'b1;
19864: pixelout<=1'b1;
19865: pixelout<=1'b1;
19866: pixelout<=1'b1;
19867: pixelout<=1'b1;
19868: pixelout<=1'b1;
19869: pixelout<=1'b1;
19870: pixelout<=1'b1;
19871: pixelout<=1'b1;
19872: pixelout<=1'b1;
19873: pixelout<=1'b1;
19874: pixelout<=1'b1;
19875: pixelout<=1'b1;
19876: pixelout<=1'b1;
19877: pixelout<=1'b1;
19878: pixelout<=1'b1;
19879: pixelout<=1'b1;
19880: pixelout<=1'b1;
19881: pixelout<=1'b1;
19882: pixelout<=1'b1;
19883: pixelout<=1'b1;
19884: pixelout<=1'b1;
19885: pixelout<=1'b1;
19886: pixelout<=1'b1;
19887: pixelout<=1'b1;
19888: pixelout<=1'b1;
19889: pixelout<=1'b1;
19890: pixelout<=1'b1;
19891: pixelout<=1'b1;
19892: pixelout<=1'b1;
19893: pixelout<=1'b1;
19894: pixelout<=1'b1;
19895: pixelout<=1'b1;
19896: pixelout<=1'b1;
19897: pixelout<=1'b1;
19898: pixelout<=1'b1;
19899: pixelout<=1'b1;
19900: pixelout<=1'b1;
19901: pixelout<=1'b1;
19902: pixelout<=1'b1;
19903: pixelout<=1'b1;
19904: pixelout<=1'b1;
19905: pixelout<=1'b1;
19906: pixelout<=1'b1;
19907: pixelout<=1'b1;
19908: pixelout<=1'b1;
19909: pixelout<=1'b1;
19910: pixelout<=1'b1;
19911: pixelout<=1'b1;
19912: pixelout<=1'b1;
19913: pixelout<=1'b1;
19914: pixelout<=1'b1;
19915: pixelout<=1'b1;
19916: pixelout<=1'b1;
19917: pixelout<=1'b1;
19918: pixelout<=1'b1;
19919: pixelout<=1'b1;
19920: pixelout<=1'b1;
19921: pixelout<=1'b1;
19922: pixelout<=1'b1;
19923: pixelout<=1'b1;
19924: pixelout<=1'b1;
19925: pixelout<=1'b1;
19926: pixelout<=1'b1;
19927: pixelout<=1'b1;
19928: pixelout<=1'b1;
19929: pixelout<=1'b1;
19930: pixelout<=1'b1;
19931: pixelout<=1'b1;
19932: pixelout<=1'b1;
19933: pixelout<=1'b1;
19934: pixelout<=1'b1;
19935: pixelout<=1'b1;
19936: pixelout<=1'b1;
19937: pixelout<=1'b1;
19938: pixelout<=1'b1;
19939: pixelout<=1'b1;
19940: pixelout<=1'b1;
19941: pixelout<=1'b1;
19942: pixelout<=1'b1;
19943: pixelout<=1'b1;
19944: pixelout<=1'b1;
19945: pixelout<=1'b1;
19946: pixelout<=1'b1;
19947: pixelout<=1'b1;
19948: pixelout<=1'b1;
19949: pixelout<=1'b1;
19950: pixelout<=1'b1;
19951: pixelout<=1'b1;
19952: pixelout<=1'b1;
19953: pixelout<=1'b1;
19954: pixelout<=1'b1;
19955: pixelout<=1'b1;
19956: pixelout<=1'b1;
19957: pixelout<=1'b1;
19958: pixelout<=1'b1;
19959: pixelout<=1'b1;
19960: pixelout<=1'b1;
19961: pixelout<=1'b1;
19962: pixelout<=1'b1;
19963: pixelout<=1'b1;
19964: pixelout<=1'b1;
19965: pixelout<=1'b1;
19966: pixelout<=1'b1;
19967: pixelout<=1'b1;
19968: pixelout<=1'b1;
19969: pixelout<=1'b1;
19970: pixelout<=1'b1;
19971: pixelout<=1'b1;
19972: pixelout<=1'b1;
19973: pixelout<=1'b1;
19974: pixelout<=1'b1;
19975: pixelout<=1'b1;
19976: pixelout<=1'b1;
19977: pixelout<=1'b1;
19978: pixelout<=1'b1;
19979: pixelout<=1'b1;
19980: pixelout<=1'b1;
19981: pixelout<=1'b1;
19982: pixelout<=1'b1;
19983: pixelout<=1'b1;
19984: pixelout<=1'b1;
19985: pixelout<=1'b1;
19986: pixelout<=1'b1;
19987: pixelout<=1'b1;
19988: pixelout<=1'b1;
19989: pixelout<=1'b1;
19990: pixelout<=1'b1;
19991: pixelout<=1'b1;
19992: pixelout<=1'b1;
19993: pixelout<=1'b1;
19994: pixelout<=1'b1;
19995: pixelout<=1'b1;
19996: pixelout<=1'b1;
19997: pixelout<=1'b1;
19998: pixelout<=1'b1;
19999: pixelout<=1'b1;
20000: pixelout<=1'b1;
20001: pixelout<=1'b1;
20002: pixelout<=1'b1;
20003: pixelout<=1'b1;
20004: pixelout<=1'b1;
20005: pixelout<=1'b1;
20006: pixelout<=1'b1;
20007: pixelout<=1'b1;
20008: pixelout<=1'b1;
20009: pixelout<=1'b1;
20010: pixelout<=1'b1;
20011: pixelout<=1'b1;
20012: pixelout<=1'b1;
20013: pixelout<=1'b1;
20014: pixelout<=1'b1;
20015: pixelout<=1'b1;
20016: pixelout<=1'b1;
20017: pixelout<=1'b1;
20018: pixelout<=1'b1;
20019: pixelout<=1'b1;
20020: pixelout<=1'b1;
20021: pixelout<=1'b1;
20022: pixelout<=1'b1;
20023: pixelout<=1'b1;
20024: pixelout<=1'b1;
20025: pixelout<=1'b1;
20026: pixelout<=1'b1;
20027: pixelout<=1'b1;
20028: pixelout<=1'b1;
20029: pixelout<=1'b1;
20030: pixelout<=1'b1;
20031: pixelout<=1'b1;
20032: pixelout<=1'b1;
20033: pixelout<=1'b1;
20034: pixelout<=1'b1;
20035: pixelout<=1'b1;
20036: pixelout<=1'b1;
20037: pixelout<=1'b1;
20038: pixelout<=1'b1;
20039: pixelout<=1'b1;
20040: pixelout<=1'b1;
20041: pixelout<=1'b1;
20042: pixelout<=1'b1;
20043: pixelout<=1'b1;
20044: pixelout<=1'b1;
20045: pixelout<=1'b1;
20046: pixelout<=1'b1;
20047: pixelout<=1'b1;
20048: pixelout<=1'b1;
20049: pixelout<=1'b1;
20050: pixelout<=1'b1;
20051: pixelout<=1'b1;
20052: pixelout<=1'b1;
20053: pixelout<=1'b1;
20054: pixelout<=1'b1;
20055: pixelout<=1'b1;
20056: pixelout<=1'b1;
20057: pixelout<=1'b1;
20058: pixelout<=1'b1;
20059: pixelout<=1'b1;
20060: pixelout<=1'b1;
20061: pixelout<=1'b1;
20062: pixelout<=1'b1;
20063: pixelout<=1'b1;
20064: pixelout<=1'b1;
20065: pixelout<=1'b1;
20066: pixelout<=1'b1;
20067: pixelout<=1'b1;
20068: pixelout<=1'b1;
20069: pixelout<=1'b1;
20070: pixelout<=1'b1;
20071: pixelout<=1'b1;
20072: pixelout<=1'b1;
20073: pixelout<=1'b1;
20074: pixelout<=1'b1;
20075: pixelout<=1'b1;
20076: pixelout<=1'b1;
20077: pixelout<=1'b1;
20078: pixelout<=1'b1;
20079: pixelout<=1'b1;
20080: pixelout<=1'b1;
20081: pixelout<=1'b1;
20082: pixelout<=1'b1;
20083: pixelout<=1'b1;
20084: pixelout<=1'b1;
20085: pixelout<=1'b1;
20086: pixelout<=1'b1;
20087: pixelout<=1'b1;
20088: pixelout<=1'b1;
20089: pixelout<=1'b1;
20090: pixelout<=1'b1;
20091: pixelout<=1'b1;
20092: pixelout<=1'b1;
20093: pixelout<=1'b1;
20094: pixelout<=1'b1;
20095: pixelout<=1'b1;
20096: pixelout<=1'b1;
20097: pixelout<=1'b1;
20098: pixelout<=1'b1;
20099: pixelout<=1'b1;
20100: pixelout<=1'b1;
20101: pixelout<=1'b1;
20102: pixelout<=1'b1;
20103: pixelout<=1'b1;
20104: pixelout<=1'b1;
20105: pixelout<=1'b1;
20106: pixelout<=1'b1;
20107: pixelout<=1'b1;
20108: pixelout<=1'b1;
20109: pixelout<=1'b1;
20110: pixelout<=1'b1;
20111: pixelout<=1'b1;
20112: pixelout<=1'b1;
20113: pixelout<=1'b1;
20114: pixelout<=1'b1;
20115: pixelout<=1'b1;
20116: pixelout<=1'b1;
20117: pixelout<=1'b1;
20118: pixelout<=1'b1;
20119: pixelout<=1'b1;
20120: pixelout<=1'b1;
20121: pixelout<=1'b1;
20122: pixelout<=1'b1;
20123: pixelout<=1'b1;
20124: pixelout<=1'b1;
20125: pixelout<=1'b1;
20126: pixelout<=1'b1;
20127: pixelout<=1'b1;
20128: pixelout<=1'b1;
20129: pixelout<=1'b1;
20130: pixelout<=1'b1;
20131: pixelout<=1'b1;
20132: pixelout<=1'b1;
20133: pixelout<=1'b1;
20134: pixelout<=1'b1;
20135: pixelout<=1'b1;
20136: pixelout<=1'b1;
20137: pixelout<=1'b1;
20138: pixelout<=1'b1;
20139: pixelout<=1'b1;
20140: pixelout<=1'b1;
20141: pixelout<=1'b1;
20142: pixelout<=1'b1;
20143: pixelout<=1'b1;
20144: pixelout<=1'b1;
20145: pixelout<=1'b1;
20146: pixelout<=1'b1;
20147: pixelout<=1'b1;
20148: pixelout<=1'b1;
20149: pixelout<=1'b1;
20150: pixelout<=1'b1;
20151: pixelout<=1'b1;
20152: pixelout<=1'b1;
20153: pixelout<=1'b1;
20154: pixelout<=1'b1;
20155: pixelout<=1'b1;
20156: pixelout<=1'b1;
20157: pixelout<=1'b1;
20158: pixelout<=1'b1;
20159: pixelout<=1'b1;
20160: pixelout<=1'b1;
20161: pixelout<=1'b1;
20162: pixelout<=1'b1;
20163: pixelout<=1'b1;
20164: pixelout<=1'b1;
20165: pixelout<=1'b1;
20166: pixelout<=1'b1;
20167: pixelout<=1'b1;
20168: pixelout<=1'b1;
20169: pixelout<=1'b1;
20170: pixelout<=1'b1;
20171: pixelout<=1'b1;
20172: pixelout<=1'b1;
20173: pixelout<=1'b1;
20174: pixelout<=1'b1;
20175: pixelout<=1'b1;
20176: pixelout<=1'b1;
20177: pixelout<=1'b1;
20178: pixelout<=1'b1;
20179: pixelout<=1'b1;
20180: pixelout<=1'b1;
20181: pixelout<=1'b1;
20182: pixelout<=1'b1;
20183: pixelout<=1'b1;
20184: pixelout<=1'b1;
20185: pixelout<=1'b1;
20186: pixelout<=1'b1;
20187: pixelout<=1'b1;
20188: pixelout<=1'b1;
20189: pixelout<=1'b1;
20190: pixelout<=1'b1;
20191: pixelout<=1'b1;
20192: pixelout<=1'b1;
20193: pixelout<=1'b1;
20194: pixelout<=1'b1;
20195: pixelout<=1'b1;
20196: pixelout<=1'b1;
20197: pixelout<=1'b1;
20198: pixelout<=1'b1;
20199: pixelout<=1'b1;
20200: pixelout<=1'b1;
20201: pixelout<=1'b1;
20202: pixelout<=1'b1;
20203: pixelout<=1'b1;
20204: pixelout<=1'b1;
20205: pixelout<=1'b1;
20206: pixelout<=1'b1;
20207: pixelout<=1'b1;
20208: pixelout<=1'b1;
20209: pixelout<=1'b1;
20210: pixelout<=1'b1;
20211: pixelout<=1'b1;
20212: pixelout<=1'b1;
20213: pixelout<=1'b1;
20214: pixelout<=1'b1;
20215: pixelout<=1'b1;
20216: pixelout<=1'b1;
20217: pixelout<=1'b1;
20218: pixelout<=1'b1;
20219: pixelout<=1'b1;
20220: pixelout<=1'b1;
20221: pixelout<=1'b1;
20222: pixelout<=1'b1;
20223: pixelout<=1'b1;
20224: pixelout<=1'b1;
20225: pixelout<=1'b1;
20226: pixelout<=1'b1;
20227: pixelout<=1'b1;
20228: pixelout<=1'b1;
20229: pixelout<=1'b1;
20230: pixelout<=1'b1;
20231: pixelout<=1'b1;
20232: pixelout<=1'b1;
20233: pixelout<=1'b1;
20234: pixelout<=1'b1;
20235: pixelout<=1'b1;
20236: pixelout<=1'b1;
20237: pixelout<=1'b1;
20238: pixelout<=1'b1;
20239: pixelout<=1'b1;
20240: pixelout<=1'b1;
20241: pixelout<=1'b1;
20242: pixelout<=1'b1;
20243: pixelout<=1'b1;
20244: pixelout<=1'b1;
20245: pixelout<=1'b1;
20246: pixelout<=1'b1;
20247: pixelout<=1'b1;
20248: pixelout<=1'b1;
20249: pixelout<=1'b1;
20250: pixelout<=1'b1;
20251: pixelout<=1'b1;
20252: pixelout<=1'b1;
20253: pixelout<=1'b1;
20254: pixelout<=1'b1;
20255: pixelout<=1'b1;
20256: pixelout<=1'b1;
20257: pixelout<=1'b1;
20258: pixelout<=1'b1;
20259: pixelout<=1'b1;
20260: pixelout<=1'b1;
20261: pixelout<=1'b1;
20262: pixelout<=1'b1;
20263: pixelout<=1'b1;
20264: pixelout<=1'b1;
20265: pixelout<=1'b1;
20266: pixelout<=1'b1;
20267: pixelout<=1'b1;
20268: pixelout<=1'b1;
20269: pixelout<=1'b1;
20270: pixelout<=1'b1;
20271: pixelout<=1'b1;
20272: pixelout<=1'b1;
20273: pixelout<=1'b1;
20274: pixelout<=1'b1;
20275: pixelout<=1'b1;
20276: pixelout<=1'b1;
20277: pixelout<=1'b1;
20278: pixelout<=1'b1;
20279: pixelout<=1'b1;
20280: pixelout<=1'b1;
20281: pixelout<=1'b1;
20282: pixelout<=1'b1;
20283: pixelout<=1'b1;
20284: pixelout<=1'b1;
20285: pixelout<=1'b1;
20286: pixelout<=1'b1;
20287: pixelout<=1'b1;
20288: pixelout<=1'b1;
20289: pixelout<=1'b1;
20290: pixelout<=1'b1;
20291: pixelout<=1'b1;
20292: pixelout<=1'b1;
20293: pixelout<=1'b1;
20294: pixelout<=1'b1;
20295: pixelout<=1'b1;
20296: pixelout<=1'b1;
20297: pixelout<=1'b1;
20298: pixelout<=1'b1;
20299: pixelout<=1'b1;
20300: pixelout<=1'b1;
20301: pixelout<=1'b1;
20302: pixelout<=1'b1;
20303: pixelout<=1'b1;
20304: pixelout<=1'b1;
20305: pixelout<=1'b1;
20306: pixelout<=1'b1;
20307: pixelout<=1'b1;
20308: pixelout<=1'b1;
20309: pixelout<=1'b1;
20310: pixelout<=1'b1;
20311: pixelout<=1'b1;
20312: pixelout<=1'b1;
20313: pixelout<=1'b1;
20314: pixelout<=1'b1;
20315: pixelout<=1'b1;
20316: pixelout<=1'b1;
20317: pixelout<=1'b1;
20318: pixelout<=1'b1;
20319: pixelout<=1'b1;
20320: pixelout<=1'b1;
20321: pixelout<=1'b1;
20322: pixelout<=1'b1;
20323: pixelout<=1'b1;
20324: pixelout<=1'b1;
20325: pixelout<=1'b1;
20326: pixelout<=1'b1;
20327: pixelout<=1'b1;
20328: pixelout<=1'b1;
20329: pixelout<=1'b1;
20330: pixelout<=1'b1;
20331: pixelout<=1'b1;
20332: pixelout<=1'b1;
20333: pixelout<=1'b1;
20334: pixelout<=1'b1;
20335: pixelout<=1'b1;
20336: pixelout<=1'b1;
20337: pixelout<=1'b1;
20338: pixelout<=1'b1;
20339: pixelout<=1'b1;
20340: pixelout<=1'b1;
20341: pixelout<=1'b1;
20342: pixelout<=1'b1;
20343: pixelout<=1'b1;
20344: pixelout<=1'b1;
20345: pixelout<=1'b1;
20346: pixelout<=1'b1;
20347: pixelout<=1'b1;
20348: pixelout<=1'b1;
20349: pixelout<=1'b1;
20350: pixelout<=1'b1;
20351: pixelout<=1'b1;
20352: pixelout<=1'b1;
20353: pixelout<=1'b1;
20354: pixelout<=1'b1;
20355: pixelout<=1'b1;
20356: pixelout<=1'b1;
20357: pixelout<=1'b1;
20358: pixelout<=1'b1;
20359: pixelout<=1'b1;
20360: pixelout<=1'b1;
20361: pixelout<=1'b1;
20362: pixelout<=1'b1;
20363: pixelout<=1'b1;
20364: pixelout<=1'b1;
20365: pixelout<=1'b1;
20366: pixelout<=1'b1;
20367: pixelout<=1'b1;
20368: pixelout<=1'b1;
20369: pixelout<=1'b1;
20370: pixelout<=1'b1;
20371: pixelout<=1'b1;
20372: pixelout<=1'b1;
20373: pixelout<=1'b1;
20374: pixelout<=1'b1;
20375: pixelout<=1'b1;
20376: pixelout<=1'b1;
20377: pixelout<=1'b1;
20378: pixelout<=1'b1;
20379: pixelout<=1'b1;
20380: pixelout<=1'b1;
20381: pixelout<=1'b1;
20382: pixelout<=1'b1;
20383: pixelout<=1'b1;
20384: pixelout<=1'b1;
20385: pixelout<=1'b1;
20386: pixelout<=1'b1;
20387: pixelout<=1'b1;
20388: pixelout<=1'b1;
20389: pixelout<=1'b1;
20390: pixelout<=1'b1;
20391: pixelout<=1'b1;
20392: pixelout<=1'b1;
20393: pixelout<=1'b1;
20394: pixelout<=1'b1;
20395: pixelout<=1'b1;
20396: pixelout<=1'b1;
20397: pixelout<=1'b1;
20398: pixelout<=1'b1;
20399: pixelout<=1'b1;
20400: pixelout<=1'b1;
20401: pixelout<=1'b1;
20402: pixelout<=1'b1;
20403: pixelout<=1'b1;
20404: pixelout<=1'b1;
20405: pixelout<=1'b1;
20406: pixelout<=1'b1;
20407: pixelout<=1'b1;
20408: pixelout<=1'b1;
20409: pixelout<=1'b1;
20410: pixelout<=1'b1;
20411: pixelout<=1'b1;
20412: pixelout<=1'b1;
20413: pixelout<=1'b1;
20414: pixelout<=1'b1;
20415: pixelout<=1'b1;
20416: pixelout<=1'b1;
20417: pixelout<=1'b1;
20418: pixelout<=1'b1;
20419: pixelout<=1'b1;
20420: pixelout<=1'b1;
20421: pixelout<=1'b1;
20422: pixelout<=1'b1;
20423: pixelout<=1'b1;
20424: pixelout<=1'b1;
20425: pixelout<=1'b1;
20426: pixelout<=1'b1;
20427: pixelout<=1'b1;
20428: pixelout<=1'b1;
20429: pixelout<=1'b1;
20430: pixelout<=1'b1;
20431: pixelout<=1'b1;
20432: pixelout<=1'b1;
20433: pixelout<=1'b1;
20434: pixelout<=1'b1;
20435: pixelout<=1'b1;
20436: pixelout<=1'b1;
20437: pixelout<=1'b1;
20438: pixelout<=1'b1;
20439: pixelout<=1'b1;
20440: pixelout<=1'b1;
20441: pixelout<=1'b1;
20442: pixelout<=1'b1;
20443: pixelout<=1'b1;
20444: pixelout<=1'b1;
20445: pixelout<=1'b1;
20446: pixelout<=1'b1;
20447: pixelout<=1'b1;
20448: pixelout<=1'b1;
20449: pixelout<=1'b1;
20450: pixelout<=1'b1;
20451: pixelout<=1'b1;
20452: pixelout<=1'b1;
20453: pixelout<=1'b1;
20454: pixelout<=1'b1;
20455: pixelout<=1'b1;
20456: pixelout<=1'b1;
20457: pixelout<=1'b1;
20458: pixelout<=1'b1;
20459: pixelout<=1'b1;
20460: pixelout<=1'b1;
20461: pixelout<=1'b1;
20462: pixelout<=1'b1;
20463: pixelout<=1'b1;
20464: pixelout<=1'b1;
20465: pixelout<=1'b1;
20466: pixelout<=1'b1;
20467: pixelout<=1'b1;
20468: pixelout<=1'b1;
20469: pixelout<=1'b1;
20470: pixelout<=1'b1;
20471: pixelout<=1'b1;
20472: pixelout<=1'b1;
20473: pixelout<=1'b1;
20474: pixelout<=1'b1;
20475: pixelout<=1'b1;
20476: pixelout<=1'b1;
20477: pixelout<=1'b1;
20478: pixelout<=1'b1;
20479: pixelout<=1'b1;
20480: pixelout<=1'b1;
20481: pixelout<=1'b1;
20482: pixelout<=1'b1;
20483: pixelout<=1'b1;
20484: pixelout<=1'b1;
20485: pixelout<=1'b1;
20486: pixelout<=1'b1;
20487: pixelout<=1'b1;
20488: pixelout<=1'b1;
20489: pixelout<=1'b1;
20490: pixelout<=1'b1;
20491: pixelout<=1'b1;
20492: pixelout<=1'b1;
20493: pixelout<=1'b1;
20494: pixelout<=1'b1;
20495: pixelout<=1'b1;
20496: pixelout<=1'b1;
20497: pixelout<=1'b1;
20498: pixelout<=1'b1;
20499: pixelout<=1'b1;
20500: pixelout<=1'b1;
20501: pixelout<=1'b1;
20502: pixelout<=1'b1;
20503: pixelout<=1'b1;
20504: pixelout<=1'b1;
20505: pixelout<=1'b1;
20506: pixelout<=1'b1;
20507: pixelout<=1'b1;
20508: pixelout<=1'b1;
20509: pixelout<=1'b1;
20510: pixelout<=1'b1;
20511: pixelout<=1'b1;
20512: pixelout<=1'b1;
20513: pixelout<=1'b1;
20514: pixelout<=1'b1;
20515: pixelout<=1'b1;
20516: pixelout<=1'b1;
20517: pixelout<=1'b1;
20518: pixelout<=1'b1;
20519: pixelout<=1'b1;
20520: pixelout<=1'b1;
20521: pixelout<=1'b1;
20522: pixelout<=1'b1;
20523: pixelout<=1'b1;
20524: pixelout<=1'b1;
20525: pixelout<=1'b1;
20526: pixelout<=1'b1;
20527: pixelout<=1'b1;
20528: pixelout<=1'b1;
20529: pixelout<=1'b1;
20530: pixelout<=1'b1;
20531: pixelout<=1'b1;
20532: pixelout<=1'b1;
20533: pixelout<=1'b1;
20534: pixelout<=1'b1;
20535: pixelout<=1'b1;
20536: pixelout<=1'b1;
20537: pixelout<=1'b1;
20538: pixelout<=1'b1;
20539: pixelout<=1'b1;
20540: pixelout<=1'b1;
20541: pixelout<=1'b1;
20542: pixelout<=1'b1;
20543: pixelout<=1'b1;
20544: pixelout<=1'b1;
20545: pixelout<=1'b1;
20546: pixelout<=1'b1;
20547: pixelout<=1'b1;
20548: pixelout<=1'b1;
20549: pixelout<=1'b1;
20550: pixelout<=1'b1;
20551: pixelout<=1'b1;
20552: pixelout<=1'b1;
20553: pixelout<=1'b1;
20554: pixelout<=1'b1;
20555: pixelout<=1'b1;
20556: pixelout<=1'b1;
20557: pixelout<=1'b1;
20558: pixelout<=1'b1;
20559: pixelout<=1'b1;
20560: pixelout<=1'b1;
20561: pixelout<=1'b1;
20562: pixelout<=1'b1;
20563: pixelout<=1'b1;
20564: pixelout<=1'b1;
20565: pixelout<=1'b1;
20566: pixelout<=1'b1;
20567: pixelout<=1'b1;
20568: pixelout<=1'b1;
20569: pixelout<=1'b1;
20570: pixelout<=1'b1;
20571: pixelout<=1'b1;
20572: pixelout<=1'b1;
20573: pixelout<=1'b1;
20574: pixelout<=1'b1;
20575: pixelout<=1'b1;
20576: pixelout<=1'b1;
20577: pixelout<=1'b1;
20578: pixelout<=1'b1;
20579: pixelout<=1'b1;
20580: pixelout<=1'b1;
20581: pixelout<=1'b1;
20582: pixelout<=1'b1;
20583: pixelout<=1'b1;
20584: pixelout<=1'b1;
20585: pixelout<=1'b1;
20586: pixelout<=1'b1;
20587: pixelout<=1'b1;
20588: pixelout<=1'b1;
20589: pixelout<=1'b1;
20590: pixelout<=1'b1;
20591: pixelout<=1'b1;
20592: pixelout<=1'b1;
20593: pixelout<=1'b1;
20594: pixelout<=1'b1;
20595: pixelout<=1'b1;
20596: pixelout<=1'b1;
20597: pixelout<=1'b1;
20598: pixelout<=1'b1;
20599: pixelout<=1'b1;
20600: pixelout<=1'b1;
20601: pixelout<=1'b1;
20602: pixelout<=1'b1;
20603: pixelout<=1'b1;
20604: pixelout<=1'b1;
20605: pixelout<=1'b1;
20606: pixelout<=1'b1;
20607: pixelout<=1'b1;
20608: pixelout<=1'b1;
20609: pixelout<=1'b1;
20610: pixelout<=1'b1;
20611: pixelout<=1'b1;
20612: pixelout<=1'b1;
20613: pixelout<=1'b1;
20614: pixelout<=1'b1;
20615: pixelout<=1'b1;
20616: pixelout<=1'b1;
20617: pixelout<=1'b1;
20618: pixelout<=1'b1;
20619: pixelout<=1'b1;
20620: pixelout<=1'b1;
20621: pixelout<=1'b1;
20622: pixelout<=1'b1;
20623: pixelout<=1'b1;
20624: pixelout<=1'b1;
20625: pixelout<=1'b1;
20626: pixelout<=1'b1;
20627: pixelout<=1'b1;
20628: pixelout<=1'b1;
20629: pixelout<=1'b1;
20630: pixelout<=1'b1;
20631: pixelout<=1'b1;
20632: pixelout<=1'b1;
20633: pixelout<=1'b1;
20634: pixelout<=1'b1;
20635: pixelout<=1'b1;
20636: pixelout<=1'b1;
20637: pixelout<=1'b1;
20638: pixelout<=1'b1;
20639: pixelout<=1'b1;
20640: pixelout<=1'b1;
20641: pixelout<=1'b1;
20642: pixelout<=1'b1;
20643: pixelout<=1'b1;
20644: pixelout<=1'b1;
20645: pixelout<=1'b1;
20646: pixelout<=1'b1;
20647: pixelout<=1'b1;
20648: pixelout<=1'b1;
20649: pixelout<=1'b1;
20650: pixelout<=1'b1;
20651: pixelout<=1'b1;
20652: pixelout<=1'b1;
20653: pixelout<=1'b1;
20654: pixelout<=1'b1;
20655: pixelout<=1'b1;
20656: pixelout<=1'b1;
20657: pixelout<=1'b1;
20658: pixelout<=1'b1;
20659: pixelout<=1'b1;
20660: pixelout<=1'b1;
20661: pixelout<=1'b1;
20662: pixelout<=1'b1;
20663: pixelout<=1'b1;
20664: pixelout<=1'b1;
20665: pixelout<=1'b1;
20666: pixelout<=1'b1;
20667: pixelout<=1'b1;
20668: pixelout<=1'b1;
20669: pixelout<=1'b1;
20670: pixelout<=1'b1;
20671: pixelout<=1'b1;
20672: pixelout<=1'b1;
20673: pixelout<=1'b1;
20674: pixelout<=1'b1;
20675: pixelout<=1'b1;
20676: pixelout<=1'b1;
20677: pixelout<=1'b1;
20678: pixelout<=1'b1;
20679: pixelout<=1'b1;
20680: pixelout<=1'b1;
20681: pixelout<=1'b1;
20682: pixelout<=1'b1;
20683: pixelout<=1'b1;
20684: pixelout<=1'b1;
20685: pixelout<=1'b1;
20686: pixelout<=1'b1;
20687: pixelout<=1'b1;
20688: pixelout<=1'b1;
20689: pixelout<=1'b1;
20690: pixelout<=1'b1;
20691: pixelout<=1'b1;
20692: pixelout<=1'b1;
20693: pixelout<=1'b1;
20694: pixelout<=1'b1;
20695: pixelout<=1'b1;
20696: pixelout<=1'b1;
20697: pixelout<=1'b1;
20698: pixelout<=1'b1;
20699: pixelout<=1'b1;
20700: pixelout<=1'b1;
20701: pixelout<=1'b1;
20702: pixelout<=1'b1;
20703: pixelout<=1'b1;
20704: pixelout<=1'b1;
20705: pixelout<=1'b1;
20706: pixelout<=1'b1;
20707: pixelout<=1'b1;
20708: pixelout<=1'b1;
20709: pixelout<=1'b1;
20710: pixelout<=1'b1;
20711: pixelout<=1'b1;
20712: pixelout<=1'b1;
20713: pixelout<=1'b1;
20714: pixelout<=1'b1;
20715: pixelout<=1'b1;
20716: pixelout<=1'b1;
20717: pixelout<=1'b1;
20718: pixelout<=1'b1;
20719: pixelout<=1'b1;
20720: pixelout<=1'b1;
20721: pixelout<=1'b1;
20722: pixelout<=1'b1;
20723: pixelout<=1'b1;
20724: pixelout<=1'b1;
20725: pixelout<=1'b1;
20726: pixelout<=1'b1;
20727: pixelout<=1'b1;
20728: pixelout<=1'b1;
20729: pixelout<=1'b1;
20730: pixelout<=1'b1;
20731: pixelout<=1'b1;
20732: pixelout<=1'b1;
20733: pixelout<=1'b1;
20734: pixelout<=1'b1;
20735: pixelout<=1'b1;
20736: pixelout<=1'b1;
20737: pixelout<=1'b1;
20738: pixelout<=1'b1;
20739: pixelout<=1'b1;
20740: pixelout<=1'b1;
20741: pixelout<=1'b1;
20742: pixelout<=1'b1;
20743: pixelout<=1'b1;
20744: pixelout<=1'b1;
20745: pixelout<=1'b1;
20746: pixelout<=1'b1;
20747: pixelout<=1'b1;
20748: pixelout<=1'b1;
20749: pixelout<=1'b1;
20750: pixelout<=1'b1;
20751: pixelout<=1'b1;
20752: pixelout<=1'b1;
20753: pixelout<=1'b1;
20754: pixelout<=1'b1;
20755: pixelout<=1'b1;
20756: pixelout<=1'b1;
20757: pixelout<=1'b1;
20758: pixelout<=1'b1;
20759: pixelout<=1'b1;
20760: pixelout<=1'b1;
20761: pixelout<=1'b1;
20762: pixelout<=1'b1;
20763: pixelout<=1'b1;
20764: pixelout<=1'b1;
20765: pixelout<=1'b1;
20766: pixelout<=1'b1;
20767: pixelout<=1'b1;
20768: pixelout<=1'b1;
20769: pixelout<=1'b1;
20770: pixelout<=1'b1;
20771: pixelout<=1'b1;
20772: pixelout<=1'b1;
20773: pixelout<=1'b1;
20774: pixelout<=1'b1;
20775: pixelout<=1'b1;
20776: pixelout<=1'b1;
20777: pixelout<=1'b1;
20778: pixelout<=1'b1;
20779: pixelout<=1'b1;
20780: pixelout<=1'b1;
20781: pixelout<=1'b1;
20782: pixelout<=1'b1;
20783: pixelout<=1'b1;
20784: pixelout<=1'b1;
20785: pixelout<=1'b1;
20786: pixelout<=1'b1;
20787: pixelout<=1'b1;
20788: pixelout<=1'b1;
20789: pixelout<=1'b1;
20790: pixelout<=1'b1;
20791: pixelout<=1'b1;
20792: pixelout<=1'b1;
20793: pixelout<=1'b1;
20794: pixelout<=1'b1;
20795: pixelout<=1'b1;
20796: pixelout<=1'b1;
20797: pixelout<=1'b1;
20798: pixelout<=1'b1;
20799: pixelout<=1'b1;
20800: pixelout<=1'b1;
20801: pixelout<=1'b1;
20802: pixelout<=1'b1;
20803: pixelout<=1'b1;
20804: pixelout<=1'b1;
20805: pixelout<=1'b1;
20806: pixelout<=1'b1;
20807: pixelout<=1'b1;
20808: pixelout<=1'b1;
20809: pixelout<=1'b1;
20810: pixelout<=1'b1;
20811: pixelout<=1'b1;
20812: pixelout<=1'b1;
20813: pixelout<=1'b1;
20814: pixelout<=1'b1;
20815: pixelout<=1'b1;
20816: pixelout<=1'b1;
20817: pixelout<=1'b1;
20818: pixelout<=1'b1;
20819: pixelout<=1'b1;
20820: pixelout<=1'b1;
20821: pixelout<=1'b1;
20822: pixelout<=1'b1;
20823: pixelout<=1'b1;
20824: pixelout<=1'b1;
20825: pixelout<=1'b1;
20826: pixelout<=1'b1;
20827: pixelout<=1'b1;
20828: pixelout<=1'b1;
20829: pixelout<=1'b1;
20830: pixelout<=1'b1;
20831: pixelout<=1'b1;
20832: pixelout<=1'b1;
20833: pixelout<=1'b1;
20834: pixelout<=1'b1;
20835: pixelout<=1'b1;
20836: pixelout<=1'b1;
20837: pixelout<=1'b1;
20838: pixelout<=1'b1;
20839: pixelout<=1'b1;
20840: pixelout<=1'b1;
20841: pixelout<=1'b1;
20842: pixelout<=1'b1;
20843: pixelout<=1'b1;
20844: pixelout<=1'b1;
20845: pixelout<=1'b1;
20846: pixelout<=1'b1;
20847: pixelout<=1'b1;
20848: pixelout<=1'b1;
20849: pixelout<=1'b1;
20850: pixelout<=1'b1;
20851: pixelout<=1'b1;
20852: pixelout<=1'b1;
20853: pixelout<=1'b1;
20854: pixelout<=1'b1;
20855: pixelout<=1'b1;
20856: pixelout<=1'b1;
20857: pixelout<=1'b1;
20858: pixelout<=1'b1;
20859: pixelout<=1'b1;
20860: pixelout<=1'b1;
20861: pixelout<=1'b1;
20862: pixelout<=1'b1;
20863: pixelout<=1'b1;
20864: pixelout<=1'b1;
20865: pixelout<=1'b1;
20866: pixelout<=1'b1;
20867: pixelout<=1'b1;
20868: pixelout<=1'b1;
20869: pixelout<=1'b1;
20870: pixelout<=1'b1;
20871: pixelout<=1'b1;
20872: pixelout<=1'b1;
20873: pixelout<=1'b1;
20874: pixelout<=1'b1;
20875: pixelout<=1'b1;
20876: pixelout<=1'b1;
20877: pixelout<=1'b1;
20878: pixelout<=1'b1;
20879: pixelout<=1'b1;
20880: pixelout<=1'b1;
20881: pixelout<=1'b1;
20882: pixelout<=1'b1;
20883: pixelout<=1'b1;
20884: pixelout<=1'b1;
20885: pixelout<=1'b1;
20886: pixelout<=1'b1;
20887: pixelout<=1'b1;
20888: pixelout<=1'b1;
20889: pixelout<=1'b1;
20890: pixelout<=1'b1;
20891: pixelout<=1'b1;
20892: pixelout<=1'b1;
20893: pixelout<=1'b1;
20894: pixelout<=1'b1;
20895: pixelout<=1'b1;
20896: pixelout<=1'b1;
20897: pixelout<=1'b1;
20898: pixelout<=1'b1;
20899: pixelout<=1'b1;
20900: pixelout<=1'b1;
20901: pixelout<=1'b1;
20902: pixelout<=1'b1;
20903: pixelout<=1'b1;
20904: pixelout<=1'b1;
20905: pixelout<=1'b1;
20906: pixelout<=1'b1;
20907: pixelout<=1'b1;
20908: pixelout<=1'b1;
20909: pixelout<=1'b1;
20910: pixelout<=1'b1;
20911: pixelout<=1'b1;
20912: pixelout<=1'b1;
20913: pixelout<=1'b1;
20914: pixelout<=1'b1;
20915: pixelout<=1'b1;
20916: pixelout<=1'b1;
20917: pixelout<=1'b1;
20918: pixelout<=1'b1;
20919: pixelout<=1'b1;
20920: pixelout<=1'b1;
20921: pixelout<=1'b1;
20922: pixelout<=1'b1;
20923: pixelout<=1'b1;
20924: pixelout<=1'b1;
20925: pixelout<=1'b1;
20926: pixelout<=1'b1;
20927: pixelout<=1'b1;
20928: pixelout<=1'b1;
20929: pixelout<=1'b1;
20930: pixelout<=1'b1;
20931: pixelout<=1'b1;
20932: pixelout<=1'b1;
20933: pixelout<=1'b1;
20934: pixelout<=1'b1;
20935: pixelout<=1'b1;
20936: pixelout<=1'b1;
20937: pixelout<=1'b1;
20938: pixelout<=1'b1;
20939: pixelout<=1'b1;
20940: pixelout<=1'b1;
20941: pixelout<=1'b1;
20942: pixelout<=1'b1;
20943: pixelout<=1'b1;
20944: pixelout<=1'b1;
20945: pixelout<=1'b1;
20946: pixelout<=1'b1;
20947: pixelout<=1'b1;
20948: pixelout<=1'b1;
20949: pixelout<=1'b1;
20950: pixelout<=1'b1;
20951: pixelout<=1'b1;
20952: pixelout<=1'b1;
20953: pixelout<=1'b1;
20954: pixelout<=1'b1;
20955: pixelout<=1'b1;
20956: pixelout<=1'b1;
20957: pixelout<=1'b1;
20958: pixelout<=1'b1;
20959: pixelout<=1'b1;
20960: pixelout<=1'b1;
20961: pixelout<=1'b1;
20962: pixelout<=1'b1;
20963: pixelout<=1'b1;
20964: pixelout<=1'b1;
20965: pixelout<=1'b1;
20966: pixelout<=1'b1;
20967: pixelout<=1'b1;
20968: pixelout<=1'b1;
20969: pixelout<=1'b1;
20970: pixelout<=1'b1;
20971: pixelout<=1'b1;
20972: pixelout<=1'b1;
20973: pixelout<=1'b1;
20974: pixelout<=1'b1;
20975: pixelout<=1'b1;
20976: pixelout<=1'b1;
20977: pixelout<=1'b1;
20978: pixelout<=1'b1;
20979: pixelout<=1'b1;
20980: pixelout<=1'b1;
20981: pixelout<=1'b1;
20982: pixelout<=1'b1;
20983: pixelout<=1'b1;
20984: pixelout<=1'b1;
20985: pixelout<=1'b1;
20986: pixelout<=1'b1;
20987: pixelout<=1'b1;
20988: pixelout<=1'b1;
20989: pixelout<=1'b1;
20990: pixelout<=1'b1;
20991: pixelout<=1'b1;
20992: pixelout<=1'b1;
20993: pixelout<=1'b1;
20994: pixelout<=1'b1;
20995: pixelout<=1'b1;
20996: pixelout<=1'b1;
20997: pixelout<=1'b1;
20998: pixelout<=1'b1;
20999: pixelout<=1'b1;
21000: pixelout<=1'b1;
21001: pixelout<=1'b1;
21002: pixelout<=1'b1;
21003: pixelout<=1'b1;
21004: pixelout<=1'b1;
21005: pixelout<=1'b1;
21006: pixelout<=1'b1;
21007: pixelout<=1'b1;
21008: pixelout<=1'b1;
21009: pixelout<=1'b1;
21010: pixelout<=1'b1;
21011: pixelout<=1'b1;
21012: pixelout<=1'b1;
21013: pixelout<=1'b1;
21014: pixelout<=1'b1;
21015: pixelout<=1'b1;
21016: pixelout<=1'b1;
21017: pixelout<=1'b1;
21018: pixelout<=1'b1;
21019: pixelout<=1'b1;
21020: pixelout<=1'b1;
21021: pixelout<=1'b1;
21022: pixelout<=1'b1;
21023: pixelout<=1'b1;
21024: pixelout<=1'b1;
21025: pixelout<=1'b1;
21026: pixelout<=1'b1;
21027: pixelout<=1'b1;
21028: pixelout<=1'b1;
21029: pixelout<=1'b1;
21030: pixelout<=1'b1;
21031: pixelout<=1'b1;
21032: pixelout<=1'b1;
21033: pixelout<=1'b1;
21034: pixelout<=1'b1;
21035: pixelout<=1'b1;
21036: pixelout<=1'b1;
21037: pixelout<=1'b1;
21038: pixelout<=1'b1;
21039: pixelout<=1'b1;
21040: pixelout<=1'b1;
21041: pixelout<=1'b1;
21042: pixelout<=1'b1;
21043: pixelout<=1'b1;
21044: pixelout<=1'b1;
21045: pixelout<=1'b1;
21046: pixelout<=1'b1;
21047: pixelout<=1'b1;
21048: pixelout<=1'b1;
21049: pixelout<=1'b1;
21050: pixelout<=1'b1;
21051: pixelout<=1'b1;
21052: pixelout<=1'b1;
21053: pixelout<=1'b1;
21054: pixelout<=1'b1;
21055: pixelout<=1'b1;
21056: pixelout<=1'b1;
21057: pixelout<=1'b1;
21058: pixelout<=1'b1;
21059: pixelout<=1'b1;
21060: pixelout<=1'b1;
21061: pixelout<=1'b1;
21062: pixelout<=1'b1;
21063: pixelout<=1'b1;
21064: pixelout<=1'b1;
21065: pixelout<=1'b1;
21066: pixelout<=1'b1;
21067: pixelout<=1'b1;
21068: pixelout<=1'b1;
21069: pixelout<=1'b1;
21070: pixelout<=1'b1;
21071: pixelout<=1'b1;
21072: pixelout<=1'b1;
21073: pixelout<=1'b1;
21074: pixelout<=1'b1;
21075: pixelout<=1'b1;
21076: pixelout<=1'b1;
21077: pixelout<=1'b1;
21078: pixelout<=1'b1;
21079: pixelout<=1'b1;
21080: pixelout<=1'b1;
21081: pixelout<=1'b1;
21082: pixelout<=1'b1;
21083: pixelout<=1'b1;
21084: pixelout<=1'b1;
21085: pixelout<=1'b1;
21086: pixelout<=1'b1;
21087: pixelout<=1'b1;
21088: pixelout<=1'b1;
21089: pixelout<=1'b1;
21090: pixelout<=1'b1;
21091: pixelout<=1'b1;
21092: pixelout<=1'b1;
21093: pixelout<=1'b1;
21094: pixelout<=1'b1;
21095: pixelout<=1'b1;
21096: pixelout<=1'b1;
21097: pixelout<=1'b1;
21098: pixelout<=1'b1;
21099: pixelout<=1'b1;
21100: pixelout<=1'b1;
21101: pixelout<=1'b1;
21102: pixelout<=1'b1;
21103: pixelout<=1'b1;
21104: pixelout<=1'b1;
21105: pixelout<=1'b1;
21106: pixelout<=1'b1;
21107: pixelout<=1'b1;
21108: pixelout<=1'b1;
21109: pixelout<=1'b1;
21110: pixelout<=1'b1;
21111: pixelout<=1'b1;
21112: pixelout<=1'b1;
21113: pixelout<=1'b1;
21114: pixelout<=1'b1;
21115: pixelout<=1'b1;
21116: pixelout<=1'b1;
21117: pixelout<=1'b1;
21118: pixelout<=1'b1;
21119: pixelout<=1'b1;
21120: pixelout<=1'b1;
21121: pixelout<=1'b1;
21122: pixelout<=1'b1;
21123: pixelout<=1'b1;
21124: pixelout<=1'b1;
21125: pixelout<=1'b1;
21126: pixelout<=1'b1;
21127: pixelout<=1'b1;
21128: pixelout<=1'b1;
21129: pixelout<=1'b1;
21130: pixelout<=1'b1;
21131: pixelout<=1'b1;
21132: pixelout<=1'b1;
21133: pixelout<=1'b1;
21134: pixelout<=1'b1;
21135: pixelout<=1'b1;
21136: pixelout<=1'b1;
21137: pixelout<=1'b1;
21138: pixelout<=1'b1;
21139: pixelout<=1'b1;
21140: pixelout<=1'b1;
21141: pixelout<=1'b1;
21142: pixelout<=1'b1;
21143: pixelout<=1'b1;
21144: pixelout<=1'b1;
21145: pixelout<=1'b1;
21146: pixelout<=1'b1;
21147: pixelout<=1'b1;
21148: pixelout<=1'b1;
21149: pixelout<=1'b1;
21150: pixelout<=1'b1;
21151: pixelout<=1'b1;
21152: pixelout<=1'b1;
21153: pixelout<=1'b1;
21154: pixelout<=1'b1;
21155: pixelout<=1'b1;
21156: pixelout<=1'b1;
21157: pixelout<=1'b1;
21158: pixelout<=1'b1;
21159: pixelout<=1'b1;
21160: pixelout<=1'b1;
21161: pixelout<=1'b1;
21162: pixelout<=1'b1;
21163: pixelout<=1'b1;
21164: pixelout<=1'b1;
21165: pixelout<=1'b1;
21166: pixelout<=1'b1;
21167: pixelout<=1'b1;
21168: pixelout<=1'b1;
21169: pixelout<=1'b1;
21170: pixelout<=1'b1;
21171: pixelout<=1'b1;
21172: pixelout<=1'b1;
21173: pixelout<=1'b1;
21174: pixelout<=1'b1;
21175: pixelout<=1'b1;
21176: pixelout<=1'b1;
21177: pixelout<=1'b1;
21178: pixelout<=1'b1;
21179: pixelout<=1'b1;
21180: pixelout<=1'b1;
21181: pixelout<=1'b1;
21182: pixelout<=1'b1;
21183: pixelout<=1'b1;
21184: pixelout<=1'b1;
21185: pixelout<=1'b1;
21186: pixelout<=1'b1;
21187: pixelout<=1'b1;
21188: pixelout<=1'b1;
21189: pixelout<=1'b1;
21190: pixelout<=1'b1;
21191: pixelout<=1'b1;
21192: pixelout<=1'b1;
21193: pixelout<=1'b1;
21194: pixelout<=1'b1;
21195: pixelout<=1'b1;
21196: pixelout<=1'b1;
21197: pixelout<=1'b1;
21198: pixelout<=1'b1;
21199: pixelout<=1'b1;
21200: pixelout<=1'b1;
21201: pixelout<=1'b1;
21202: pixelout<=1'b1;
21203: pixelout<=1'b1;
21204: pixelout<=1'b1;
21205: pixelout<=1'b1;
21206: pixelout<=1'b1;
21207: pixelout<=1'b1;
21208: pixelout<=1'b1;
21209: pixelout<=1'b1;
21210: pixelout<=1'b1;
21211: pixelout<=1'b1;
21212: pixelout<=1'b1;
21213: pixelout<=1'b1;
21214: pixelout<=1'b1;
21215: pixelout<=1'b1;
21216: pixelout<=1'b1;
21217: pixelout<=1'b1;
21218: pixelout<=1'b1;
21219: pixelout<=1'b1;
21220: pixelout<=1'b1;
21221: pixelout<=1'b1;
21222: pixelout<=1'b1;
21223: pixelout<=1'b1;
21224: pixelout<=1'b1;
21225: pixelout<=1'b1;
21226: pixelout<=1'b1;
21227: pixelout<=1'b1;
21228: pixelout<=1'b1;
21229: pixelout<=1'b1;
21230: pixelout<=1'b1;
21231: pixelout<=1'b1;
21232: pixelout<=1'b1;
21233: pixelout<=1'b1;
21234: pixelout<=1'b1;
21235: pixelout<=1'b1;
21236: pixelout<=1'b1;
21237: pixelout<=1'b1;
21238: pixelout<=1'b1;
21239: pixelout<=1'b1;
21240: pixelout<=1'b1;
21241: pixelout<=1'b1;
21242: pixelout<=1'b1;
21243: pixelout<=1'b1;
21244: pixelout<=1'b1;
21245: pixelout<=1'b1;
21246: pixelout<=1'b1;
21247: pixelout<=1'b1;
21248: pixelout<=1'b1;
21249: pixelout<=1'b1;
21250: pixelout<=1'b1;
21251: pixelout<=1'b1;
21252: pixelout<=1'b1;
21253: pixelout<=1'b1;
21254: pixelout<=1'b1;
21255: pixelout<=1'b1;
21256: pixelout<=1'b1;
21257: pixelout<=1'b1;
21258: pixelout<=1'b1;
21259: pixelout<=1'b1;
21260: pixelout<=1'b1;
21261: pixelout<=1'b1;
21262: pixelout<=1'b1;
21263: pixelout<=1'b1;
21264: pixelout<=1'b1;
21265: pixelout<=1'b1;
21266: pixelout<=1'b1;
21267: pixelout<=1'b1;
21268: pixelout<=1'b1;
21269: pixelout<=1'b1;
21270: pixelout<=1'b1;
21271: pixelout<=1'b1;
21272: pixelout<=1'b1;
21273: pixelout<=1'b1;
21274: pixelout<=1'b1;
21275: pixelout<=1'b1;
21276: pixelout<=1'b1;
21277: pixelout<=1'b1;
21278: pixelout<=1'b1;
21279: pixelout<=1'b1;
21280: pixelout<=1'b1;
21281: pixelout<=1'b1;
21282: pixelout<=1'b1;
21283: pixelout<=1'b1;
21284: pixelout<=1'b1;
21285: pixelout<=1'b1;
21286: pixelout<=1'b1;
21287: pixelout<=1'b1;
21288: pixelout<=1'b1;
21289: pixelout<=1'b1;
21290: pixelout<=1'b1;
21291: pixelout<=1'b1;
21292: pixelout<=1'b1;
21293: pixelout<=1'b1;
21294: pixelout<=1'b1;
21295: pixelout<=1'b1;
21296: pixelout<=1'b1;
21297: pixelout<=1'b1;
21298: pixelout<=1'b1;
21299: pixelout<=1'b1;
21300: pixelout<=1'b1;
21301: pixelout<=1'b1;
21302: pixelout<=1'b1;
21303: pixelout<=1'b1;
21304: pixelout<=1'b1;
21305: pixelout<=1'b1;
21306: pixelout<=1'b1;
21307: pixelout<=1'b1;
21308: pixelout<=1'b1;
21309: pixelout<=1'b1;
21310: pixelout<=1'b1;
21311: pixelout<=1'b1;
21312: pixelout<=1'b1;
21313: pixelout<=1'b1;
21314: pixelout<=1'b1;
21315: pixelout<=1'b1;
21316: pixelout<=1'b1;
21317: pixelout<=1'b1;
21318: pixelout<=1'b1;
21319: pixelout<=1'b1;
21320: pixelout<=1'b1;
21321: pixelout<=1'b1;
21322: pixelout<=1'b1;
21323: pixelout<=1'b1;
21324: pixelout<=1'b1;
21325: pixelout<=1'b1;
21326: pixelout<=1'b1;
21327: pixelout<=1'b1;
21328: pixelout<=1'b1;
21329: pixelout<=1'b1;
21330: pixelout<=1'b1;
21331: pixelout<=1'b1;
21332: pixelout<=1'b1;
21333: pixelout<=1'b1;
21334: pixelout<=1'b1;
21335: pixelout<=1'b1;
21336: pixelout<=1'b1;
21337: pixelout<=1'b1;
21338: pixelout<=1'b1;
21339: pixelout<=1'b1;
21340: pixelout<=1'b1;
21341: pixelout<=1'b1;
21342: pixelout<=1'b1;
21343: pixelout<=1'b1;
21344: pixelout<=1'b1;
21345: pixelout<=1'b1;
21346: pixelout<=1'b1;
21347: pixelout<=1'b1;
21348: pixelout<=1'b1;
21349: pixelout<=1'b1;
21350: pixelout<=1'b1;
21351: pixelout<=1'b1;
21352: pixelout<=1'b1;
21353: pixelout<=1'b1;
21354: pixelout<=1'b1;
21355: pixelout<=1'b1;
21356: pixelout<=1'b1;
21357: pixelout<=1'b1;
21358: pixelout<=1'b1;
21359: pixelout<=1'b1;
21360: pixelout<=1'b1;
21361: pixelout<=1'b1;
21362: pixelout<=1'b1;
21363: pixelout<=1'b1;
21364: pixelout<=1'b1;
21365: pixelout<=1'b1;
21366: pixelout<=1'b1;
21367: pixelout<=1'b1;
21368: pixelout<=1'b1;
21369: pixelout<=1'b1;
21370: pixelout<=1'b1;
21371: pixelout<=1'b1;
21372: pixelout<=1'b1;
21373: pixelout<=1'b1;
21374: pixelout<=1'b1;
21375: pixelout<=1'b1;
21376: pixelout<=1'b1;
21377: pixelout<=1'b1;
21378: pixelout<=1'b1;
21379: pixelout<=1'b1;
21380: pixelout<=1'b1;
21381: pixelout<=1'b1;
21382: pixelout<=1'b1;
21383: pixelout<=1'b1;
21384: pixelout<=1'b1;
21385: pixelout<=1'b1;
21386: pixelout<=1'b1;
21387: pixelout<=1'b1;
21388: pixelout<=1'b1;
21389: pixelout<=1'b1;
21390: pixelout<=1'b1;
21391: pixelout<=1'b1;
21392: pixelout<=1'b1;
21393: pixelout<=1'b1;
21394: pixelout<=1'b1;
21395: pixelout<=1'b1;
21396: pixelout<=1'b1;
21397: pixelout<=1'b1;
21398: pixelout<=1'b1;
21399: pixelout<=1'b1;
21400: pixelout<=1'b1;
21401: pixelout<=1'b1;
21402: pixelout<=1'b1;
21403: pixelout<=1'b1;
21404: pixelout<=1'b1;
21405: pixelout<=1'b1;
21406: pixelout<=1'b1;
21407: pixelout<=1'b1;
21408: pixelout<=1'b1;
21409: pixelout<=1'b1;
21410: pixelout<=1'b1;
21411: pixelout<=1'b1;
21412: pixelout<=1'b1;
21413: pixelout<=1'b1;
21414: pixelout<=1'b1;
21415: pixelout<=1'b1;
21416: pixelout<=1'b1;
21417: pixelout<=1'b1;
21418: pixelout<=1'b1;
21419: pixelout<=1'b1;
21420: pixelout<=1'b1;
21421: pixelout<=1'b1;
21422: pixelout<=1'b1;
21423: pixelout<=1'b1;
21424: pixelout<=1'b1;
21425: pixelout<=1'b1;
21426: pixelout<=1'b1;
21427: pixelout<=1'b1;
21428: pixelout<=1'b1;
21429: pixelout<=1'b1;
21430: pixelout<=1'b1;
21431: pixelout<=1'b1;
21432: pixelout<=1'b1;
21433: pixelout<=1'b1;
21434: pixelout<=1'b1;
21435: pixelout<=1'b1;
21436: pixelout<=1'b1;
21437: pixelout<=1'b1;
21438: pixelout<=1'b1;
21439: pixelout<=1'b1;
21440: pixelout<=1'b1;
21441: pixelout<=1'b1;
21442: pixelout<=1'b1;
21443: pixelout<=1'b1;
21444: pixelout<=1'b1;
21445: pixelout<=1'b1;
21446: pixelout<=1'b1;
21447: pixelout<=1'b1;
21448: pixelout<=1'b1;
21449: pixelout<=1'b1;
21450: pixelout<=1'b1;
21451: pixelout<=1'b1;
21452: pixelout<=1'b1;
21453: pixelout<=1'b1;
21454: pixelout<=1'b1;
21455: pixelout<=1'b1;
21456: pixelout<=1'b1;
21457: pixelout<=1'b1;
21458: pixelout<=1'b1;
21459: pixelout<=1'b1;
21460: pixelout<=1'b1;
21461: pixelout<=1'b1;
21462: pixelout<=1'b1;
21463: pixelout<=1'b1;
21464: pixelout<=1'b1;
21465: pixelout<=1'b1;
21466: pixelout<=1'b1;
21467: pixelout<=1'b1;
21468: pixelout<=1'b1;
21469: pixelout<=1'b1;
21470: pixelout<=1'b1;
21471: pixelout<=1'b1;
21472: pixelout<=1'b1;
21473: pixelout<=1'b1;
21474: pixelout<=1'b1;
21475: pixelout<=1'b1;
21476: pixelout<=1'b1;
21477: pixelout<=1'b1;
21478: pixelout<=1'b1;
21479: pixelout<=1'b1;
21480: pixelout<=1'b1;
21481: pixelout<=1'b1;
21482: pixelout<=1'b1;
21483: pixelout<=1'b1;
21484: pixelout<=1'b1;
21485: pixelout<=1'b1;
21486: pixelout<=1'b1;
21487: pixelout<=1'b1;
21488: pixelout<=1'b1;
21489: pixelout<=1'b1;
21490: pixelout<=1'b1;
21491: pixelout<=1'b1;
21492: pixelout<=1'b1;
21493: pixelout<=1'b1;
21494: pixelout<=1'b1;
21495: pixelout<=1'b1;
21496: pixelout<=1'b1;
21497: pixelout<=1'b1;
21498: pixelout<=1'b1;
21499: pixelout<=1'b1;
21500: pixelout<=1'b1;
21501: pixelout<=1'b0;
21502: pixelout<=1'b1;
21503: pixelout<=1'b1;
21504: pixelout<=1'b1;
21505: pixelout<=1'b1;
21506: pixelout<=1'b1;
21507: pixelout<=1'b1;
21508: pixelout<=1'b1;
21509: pixelout<=1'b1;
21510: pixelout<=1'b1;
21511: pixelout<=1'b1;
21512: pixelout<=1'b1;
21513: pixelout<=1'b1;
21514: pixelout<=1'b1;
21515: pixelout<=1'b1;
21516: pixelout<=1'b1;
21517: pixelout<=1'b1;
21518: pixelout<=1'b1;
21519: pixelout<=1'b1;
21520: pixelout<=1'b1;
21521: pixelout<=1'b1;
21522: pixelout<=1'b1;
21523: pixelout<=1'b1;
21524: pixelout<=1'b1;
21525: pixelout<=1'b1;
21526: pixelout<=1'b1;
21527: pixelout<=1'b1;
21528: pixelout<=1'b1;
21529: pixelout<=1'b1;
21530: pixelout<=1'b1;
21531: pixelout<=1'b1;
21532: pixelout<=1'b1;
21533: pixelout<=1'b1;
21534: pixelout<=1'b1;
21535: pixelout<=1'b1;
21536: pixelout<=1'b1;
21537: pixelout<=1'b1;
21538: pixelout<=1'b1;
21539: pixelout<=1'b1;
21540: pixelout<=1'b1;
21541: pixelout<=1'b1;
21542: pixelout<=1'b1;
21543: pixelout<=1'b1;
21544: pixelout<=1'b1;
21545: pixelout<=1'b1;
21546: pixelout<=1'b1;
21547: pixelout<=1'b1;
21548: pixelout<=1'b1;
21549: pixelout<=1'b1;
21550: pixelout<=1'b1;
21551: pixelout<=1'b1;
21552: pixelout<=1'b1;
21553: pixelout<=1'b1;
21554: pixelout<=1'b1;
21555: pixelout<=1'b1;
21556: pixelout<=1'b1;
21557: pixelout<=1'b1;
21558: pixelout<=1'b1;
21559: pixelout<=1'b1;
21560: pixelout<=1'b1;
21561: pixelout<=1'b1;
21562: pixelout<=1'b1;
21563: pixelout<=1'b1;
21564: pixelout<=1'b1;
21565: pixelout<=1'b1;
21566: pixelout<=1'b1;
21567: pixelout<=1'b1;
21568: pixelout<=1'b1;
21569: pixelout<=1'b1;
21570: pixelout<=1'b1;
21571: pixelout<=1'b1;
21572: pixelout<=1'b1;
21573: pixelout<=1'b1;
21574: pixelout<=1'b1;
21575: pixelout<=1'b1;
21576: pixelout<=1'b1;
21577: pixelout<=1'b1;
21578: pixelout<=1'b1;
21579: pixelout<=1'b1;
21580: pixelout<=1'b1;
21581: pixelout<=1'b1;
21582: pixelout<=1'b1;
21583: pixelout<=1'b1;
21584: pixelout<=1'b1;
21585: pixelout<=1'b1;
21586: pixelout<=1'b1;
21587: pixelout<=1'b1;
21588: pixelout<=1'b1;
21589: pixelout<=1'b1;
21590: pixelout<=1'b1;
21591: pixelout<=1'b1;
21592: pixelout<=1'b1;
21593: pixelout<=1'b1;
21594: pixelout<=1'b1;
21595: pixelout<=1'b1;
21596: pixelout<=1'b1;
21597: pixelout<=1'b1;
21598: pixelout<=1'b1;
21599: pixelout<=1'b1;
21600: pixelout<=1'b1;
21601: pixelout<=1'b1;
21602: pixelout<=1'b1;
21603: pixelout<=1'b1;
21604: pixelout<=1'b1;
21605: pixelout<=1'b1;
21606: pixelout<=1'b1;
21607: pixelout<=1'b1;
21608: pixelout<=1'b1;
21609: pixelout<=1'b1;
21610: pixelout<=1'b1;
21611: pixelout<=1'b1;
21612: pixelout<=1'b1;
21613: pixelout<=1'b1;
21614: pixelout<=1'b1;
21615: pixelout<=1'b1;
21616: pixelout<=1'b1;
21617: pixelout<=1'b1;
21618: pixelout<=1'b1;
21619: pixelout<=1'b1;
21620: pixelout<=1'b1;
21621: pixelout<=1'b1;
21622: pixelout<=1'b1;
21623: pixelout<=1'b1;
21624: pixelout<=1'b1;
21625: pixelout<=1'b1;
21626: pixelout<=1'b1;
21627: pixelout<=1'b1;
21628: pixelout<=1'b1;
21629: pixelout<=1'b1;
21630: pixelout<=1'b1;
21631: pixelout<=1'b1;
21632: pixelout<=1'b1;
21633: pixelout<=1'b1;
21634: pixelout<=1'b1;
21635: pixelout<=1'b1;
21636: pixelout<=1'b1;
21637: pixelout<=1'b1;
21638: pixelout<=1'b1;
21639: pixelout<=1'b1;
21640: pixelout<=1'b1;
21641: pixelout<=1'b1;
21642: pixelout<=1'b1;
21643: pixelout<=1'b1;
21644: pixelout<=1'b1;
21645: pixelout<=1'b1;
21646: pixelout<=1'b1;
21647: pixelout<=1'b1;
21648: pixelout<=1'b1;
21649: pixelout<=1'b1;
21650: pixelout<=1'b1;
21651: pixelout<=1'b1;
21652: pixelout<=1'b1;
21653: pixelout<=1'b1;
21654: pixelout<=1'b1;
21655: pixelout<=1'b1;
21656: pixelout<=1'b1;
21657: pixelout<=1'b1;
21658: pixelout<=1'b1;
21659: pixelout<=1'b1;
21660: pixelout<=1'b1;
21661: pixelout<=1'b1;
21662: pixelout<=1'b1;
21663: pixelout<=1'b1;
21664: pixelout<=1'b1;
21665: pixelout<=1'b1;
21666: pixelout<=1'b1;
21667: pixelout<=1'b1;
21668: pixelout<=1'b1;
21669: pixelout<=1'b1;
21670: pixelout<=1'b1;
21671: pixelout<=1'b1;
21672: pixelout<=1'b1;
21673: pixelout<=1'b1;
21674: pixelout<=1'b1;
21675: pixelout<=1'b1;
21676: pixelout<=1'b1;
21677: pixelout<=1'b1;
21678: pixelout<=1'b1;
21679: pixelout<=1'b1;
21680: pixelout<=1'b1;
21681: pixelout<=1'b1;
21682: pixelout<=1'b1;
21683: pixelout<=1'b1;
21684: pixelout<=1'b1;
21685: pixelout<=1'b1;
21686: pixelout<=1'b1;
21687: pixelout<=1'b1;
21688: pixelout<=1'b1;
21689: pixelout<=1'b1;
21690: pixelout<=1'b1;
21691: pixelout<=1'b1;
21692: pixelout<=1'b1;
21693: pixelout<=1'b1;
21694: pixelout<=1'b1;
21695: pixelout<=1'b1;
21696: pixelout<=1'b1;
21697: pixelout<=1'b1;
21698: pixelout<=1'b1;
21699: pixelout<=1'b1;
21700: pixelout<=1'b1;
21701: pixelout<=1'b1;
21702: pixelout<=1'b1;
21703: pixelout<=1'b1;
21704: pixelout<=1'b1;
21705: pixelout<=1'b1;
21706: pixelout<=1'b1;
21707: pixelout<=1'b1;
21708: pixelout<=1'b1;
21709: pixelout<=1'b1;
21710: pixelout<=1'b1;
21711: pixelout<=1'b1;
21712: pixelout<=1'b1;
21713: pixelout<=1'b1;
21714: pixelout<=1'b1;
21715: pixelout<=1'b1;
21716: pixelout<=1'b1;
21717: pixelout<=1'b1;
21718: pixelout<=1'b1;
21719: pixelout<=1'b1;
21720: pixelout<=1'b1;
21721: pixelout<=1'b1;
21722: pixelout<=1'b1;
21723: pixelout<=1'b0;
21724: pixelout<=1'b0;
21725: pixelout<=1'b0;
21726: pixelout<=1'b1;
21727: pixelout<=1'b1;
21728: pixelout<=1'b1;
21729: pixelout<=1'b1;
21730: pixelout<=1'b0;
21731: pixelout<=1'b0;
21732: pixelout<=1'b1;
21733: pixelout<=1'b1;
21734: pixelout<=1'b1;
21735: pixelout<=1'b0;
21736: pixelout<=1'b0;
21737: pixelout<=1'b0;
21738: pixelout<=1'b0;
21739: pixelout<=1'b1;
21740: pixelout<=1'b1;
21741: pixelout<=1'b0;
21742: pixelout<=1'b1;
21743: pixelout<=1'b1;
21744: pixelout<=1'b1;
21745: pixelout<=1'b1;
21746: pixelout<=1'b1;
21747: pixelout<=1'b1;
21748: pixelout<=1'b1;
21749: pixelout<=1'b1;
21750: pixelout<=1'b1;
21751: pixelout<=1'b1;
21752: pixelout<=1'b1;
21753: pixelout<=1'b1;
21754: pixelout<=1'b1;
21755: pixelout<=1'b1;
21756: pixelout<=1'b1;
21757: pixelout<=1'b1;
21758: pixelout<=1'b1;
21759: pixelout<=1'b1;
21760: pixelout<=1'b1;
21761: pixelout<=1'b1;
21762: pixelout<=1'b1;
21763: pixelout<=1'b1;
21764: pixelout<=1'b1;
21765: pixelout<=1'b1;
21766: pixelout<=1'b1;
21767: pixelout<=1'b1;
21768: pixelout<=1'b1;
21769: pixelout<=1'b1;
21770: pixelout<=1'b1;
21771: pixelout<=1'b1;
21772: pixelout<=1'b1;
21773: pixelout<=1'b1;
21774: pixelout<=1'b1;
21775: pixelout<=1'b1;
21776: pixelout<=1'b1;
21777: pixelout<=1'b1;
21778: pixelout<=1'b1;
21779: pixelout<=1'b1;
21780: pixelout<=1'b1;
21781: pixelout<=1'b1;
21782: pixelout<=1'b1;
21783: pixelout<=1'b1;
21784: pixelout<=1'b1;
21785: pixelout<=1'b1;
21786: pixelout<=1'b1;
21787: pixelout<=1'b1;
21788: pixelout<=1'b1;
21789: pixelout<=1'b1;
21790: pixelout<=1'b1;
21791: pixelout<=1'b1;
21792: pixelout<=1'b1;
21793: pixelout<=1'b1;
21794: pixelout<=1'b1;
21795: pixelout<=1'b1;
21796: pixelout<=1'b1;
21797: pixelout<=1'b1;
21798: pixelout<=1'b1;
21799: pixelout<=1'b1;
21800: pixelout<=1'b1;
21801: pixelout<=1'b1;
21802: pixelout<=1'b1;
21803: pixelout<=1'b1;
21804: pixelout<=1'b1;
21805: pixelout<=1'b1;
21806: pixelout<=1'b1;
21807: pixelout<=1'b1;
21808: pixelout<=1'b1;
21809: pixelout<=1'b1;
21810: pixelout<=1'b1;
21811: pixelout<=1'b1;
21812: pixelout<=1'b1;
21813: pixelout<=1'b1;
21814: pixelout<=1'b1;
21815: pixelout<=1'b1;
21816: pixelout<=1'b1;
21817: pixelout<=1'b1;
21818: pixelout<=1'b1;
21819: pixelout<=1'b1;
21820: pixelout<=1'b1;
21821: pixelout<=1'b1;
21822: pixelout<=1'b1;
21823: pixelout<=1'b1;
21824: pixelout<=1'b1;
21825: pixelout<=1'b1;
21826: pixelout<=1'b1;
21827: pixelout<=1'b1;
21828: pixelout<=1'b1;
21829: pixelout<=1'b1;
21830: pixelout<=1'b1;
21831: pixelout<=1'b1;
21832: pixelout<=1'b1;
21833: pixelout<=1'b1;
21834: pixelout<=1'b1;
21835: pixelout<=1'b1;
21836: pixelout<=1'b1;
21837: pixelout<=1'b1;
21838: pixelout<=1'b1;
21839: pixelout<=1'b1;
21840: pixelout<=1'b1;
21841: pixelout<=1'b1;
21842: pixelout<=1'b1;
21843: pixelout<=1'b1;
21844: pixelout<=1'b1;
21845: pixelout<=1'b1;
21846: pixelout<=1'b1;
21847: pixelout<=1'b1;
21848: pixelout<=1'b1;
21849: pixelout<=1'b1;
21850: pixelout<=1'b1;
21851: pixelout<=1'b1;
21852: pixelout<=1'b1;
21853: pixelout<=1'b1;
21854: pixelout<=1'b1;
21855: pixelout<=1'b1;
21856: pixelout<=1'b1;
21857: pixelout<=1'b1;
21858: pixelout<=1'b1;
21859: pixelout<=1'b1;
21860: pixelout<=1'b1;
21861: pixelout<=1'b1;
21862: pixelout<=1'b1;
21863: pixelout<=1'b1;
21864: pixelout<=1'b1;
21865: pixelout<=1'b1;
21866: pixelout<=1'b1;
21867: pixelout<=1'b1;
21868: pixelout<=1'b1;
21869: pixelout<=1'b1;
21870: pixelout<=1'b1;
21871: pixelout<=1'b1;
21872: pixelout<=1'b1;
21873: pixelout<=1'b1;
21874: pixelout<=1'b1;
21875: pixelout<=1'b1;
21876: pixelout<=1'b1;
21877: pixelout<=1'b1;
21878: pixelout<=1'b1;
21879: pixelout<=1'b1;
21880: pixelout<=1'b1;
21881: pixelout<=1'b1;
21882: pixelout<=1'b1;
21883: pixelout<=1'b1;
21884: pixelout<=1'b1;
21885: pixelout<=1'b1;
21886: pixelout<=1'b1;
21887: pixelout<=1'b1;
21888: pixelout<=1'b1;
21889: pixelout<=1'b1;
21890: pixelout<=1'b1;
21891: pixelout<=1'b1;
21892: pixelout<=1'b1;
21893: pixelout<=1'b1;
21894: pixelout<=1'b1;
21895: pixelout<=1'b1;
21896: pixelout<=1'b1;
21897: pixelout<=1'b1;
21898: pixelout<=1'b1;
21899: pixelout<=1'b1;
21900: pixelout<=1'b1;
21901: pixelout<=1'b1;
21902: pixelout<=1'b1;
21903: pixelout<=1'b1;
21904: pixelout<=1'b1;
21905: pixelout<=1'b1;
21906: pixelout<=1'b1;
21907: pixelout<=1'b1;
21908: pixelout<=1'b1;
21909: pixelout<=1'b1;
21910: pixelout<=1'b1;
21911: pixelout<=1'b1;
21912: pixelout<=1'b1;
21913: pixelout<=1'b1;
21914: pixelout<=1'b1;
21915: pixelout<=1'b1;
21916: pixelout<=1'b1;
21917: pixelout<=1'b1;
21918: pixelout<=1'b1;
21919: pixelout<=1'b1;
21920: pixelout<=1'b1;
21921: pixelout<=1'b1;
21922: pixelout<=1'b1;
21923: pixelout<=1'b1;
21924: pixelout<=1'b1;
21925: pixelout<=1'b1;
21926: pixelout<=1'b1;
21927: pixelout<=1'b1;
21928: pixelout<=1'b1;
21929: pixelout<=1'b1;
21930: pixelout<=1'b1;
21931: pixelout<=1'b1;
21932: pixelout<=1'b1;
21933: pixelout<=1'b1;
21934: pixelout<=1'b1;
21935: pixelout<=1'b1;
21936: pixelout<=1'b1;
21937: pixelout<=1'b1;
21938: pixelout<=1'b1;
21939: pixelout<=1'b1;
21940: pixelout<=1'b1;
21941: pixelout<=1'b1;
21942: pixelout<=1'b1;
21943: pixelout<=1'b1;
21944: pixelout<=1'b1;
21945: pixelout<=1'b1;
21946: pixelout<=1'b1;
21947: pixelout<=1'b1;
21948: pixelout<=1'b1;
21949: pixelout<=1'b1;
21950: pixelout<=1'b1;
21951: pixelout<=1'b1;
21952: pixelout<=1'b1;
21953: pixelout<=1'b1;
21954: pixelout<=1'b1;
21955: pixelout<=1'b1;
21956: pixelout<=1'b1;
21957: pixelout<=1'b1;
21958: pixelout<=1'b1;
21959: pixelout<=1'b1;
21960: pixelout<=1'b1;
21961: pixelout<=1'b1;
21962: pixelout<=1'b0;
21963: pixelout<=1'b1;
21964: pixelout<=1'b1;
21965: pixelout<=1'b1;
21966: pixelout<=1'b0;
21967: pixelout<=1'b1;
21968: pixelout<=1'b0;
21969: pixelout<=1'b1;
21970: pixelout<=1'b1;
21971: pixelout<=1'b1;
21972: pixelout<=1'b1;
21973: pixelout<=1'b1;
21974: pixelout<=1'b1;
21975: pixelout<=1'b1;
21976: pixelout<=1'b1;
21977: pixelout<=1'b1;
21978: pixelout<=1'b1;
21979: pixelout<=1'b1;
21980: pixelout<=1'b1;
21981: pixelout<=1'b0;
21982: pixelout<=1'b1;
21983: pixelout<=1'b1;
21984: pixelout<=1'b1;
21985: pixelout<=1'b1;
21986: pixelout<=1'b1;
21987: pixelout<=1'b1;
21988: pixelout<=1'b1;
21989: pixelout<=1'b1;
21990: pixelout<=1'b1;
21991: pixelout<=1'b1;
21992: pixelout<=1'b1;
21993: pixelout<=1'b1;
21994: pixelout<=1'b1;
21995: pixelout<=1'b1;
21996: pixelout<=1'b1;
21997: pixelout<=1'b1;
21998: pixelout<=1'b1;
21999: pixelout<=1'b1;
22000: pixelout<=1'b1;
22001: pixelout<=1'b1;
22002: pixelout<=1'b1;
22003: pixelout<=1'b1;
22004: pixelout<=1'b1;
22005: pixelout<=1'b1;
22006: pixelout<=1'b1;
22007: pixelout<=1'b1;
22008: pixelout<=1'b1;
22009: pixelout<=1'b1;
22010: pixelout<=1'b1;
22011: pixelout<=1'b1;
22012: pixelout<=1'b1;
22013: pixelout<=1'b1;
22014: pixelout<=1'b1;
22015: pixelout<=1'b1;
22016: pixelout<=1'b1;
22017: pixelout<=1'b1;
22018: pixelout<=1'b1;
22019: pixelout<=1'b1;
22020: pixelout<=1'b1;
22021: pixelout<=1'b1;
22022: pixelout<=1'b1;
22023: pixelout<=1'b1;
22024: pixelout<=1'b1;
22025: pixelout<=1'b1;
22026: pixelout<=1'b1;
22027: pixelout<=1'b1;
22028: pixelout<=1'b1;
22029: pixelout<=1'b1;
22030: pixelout<=1'b1;
22031: pixelout<=1'b1;
22032: pixelout<=1'b1;
22033: pixelout<=1'b1;
22034: pixelout<=1'b1;
22035: pixelout<=1'b1;
22036: pixelout<=1'b1;
22037: pixelout<=1'b1;
22038: pixelout<=1'b1;
22039: pixelout<=1'b1;
22040: pixelout<=1'b1;
22041: pixelout<=1'b1;
22042: pixelout<=1'b1;
22043: pixelout<=1'b1;
22044: pixelout<=1'b1;
22045: pixelout<=1'b1;
22046: pixelout<=1'b1;
22047: pixelout<=1'b1;
22048: pixelout<=1'b1;
22049: pixelout<=1'b1;
22050: pixelout<=1'b1;
22051: pixelout<=1'b1;
22052: pixelout<=1'b1;
22053: pixelout<=1'b1;
22054: pixelout<=1'b1;
22055: pixelout<=1'b1;
22056: pixelout<=1'b1;
22057: pixelout<=1'b1;
22058: pixelout<=1'b1;
22059: pixelout<=1'b1;
22060: pixelout<=1'b1;
22061: pixelout<=1'b1;
22062: pixelout<=1'b1;
22063: pixelout<=1'b1;
22064: pixelout<=1'b1;
22065: pixelout<=1'b1;
22066: pixelout<=1'b1;
22067: pixelout<=1'b1;
22068: pixelout<=1'b1;
22069: pixelout<=1'b1;
22070: pixelout<=1'b1;
22071: pixelout<=1'b1;
22072: pixelout<=1'b1;
22073: pixelout<=1'b1;
22074: pixelout<=1'b1;
22075: pixelout<=1'b1;
22076: pixelout<=1'b1;
22077: pixelout<=1'b1;
22078: pixelout<=1'b1;
22079: pixelout<=1'b1;
22080: pixelout<=1'b1;
22081: pixelout<=1'b1;
22082: pixelout<=1'b1;
22083: pixelout<=1'b1;
22084: pixelout<=1'b1;
22085: pixelout<=1'b1;
22086: pixelout<=1'b1;
22087: pixelout<=1'b1;
22088: pixelout<=1'b1;
22089: pixelout<=1'b1;
22090: pixelout<=1'b1;
22091: pixelout<=1'b1;
22092: pixelout<=1'b1;
22093: pixelout<=1'b1;
22094: pixelout<=1'b1;
22095: pixelout<=1'b1;
22096: pixelout<=1'b1;
22097: pixelout<=1'b1;
22098: pixelout<=1'b1;
22099: pixelout<=1'b1;
22100: pixelout<=1'b1;
22101: pixelout<=1'b1;
22102: pixelout<=1'b1;
22103: pixelout<=1'b1;
22104: pixelout<=1'b1;
22105: pixelout<=1'b1;
22106: pixelout<=1'b1;
22107: pixelout<=1'b1;
22108: pixelout<=1'b1;
22109: pixelout<=1'b1;
22110: pixelout<=1'b1;
22111: pixelout<=1'b1;
22112: pixelout<=1'b1;
22113: pixelout<=1'b1;
22114: pixelout<=1'b1;
22115: pixelout<=1'b1;
22116: pixelout<=1'b1;
22117: pixelout<=1'b1;
22118: pixelout<=1'b1;
22119: pixelout<=1'b1;
22120: pixelout<=1'b1;
22121: pixelout<=1'b1;
22122: pixelout<=1'b1;
22123: pixelout<=1'b1;
22124: pixelout<=1'b1;
22125: pixelout<=1'b1;
22126: pixelout<=1'b1;
22127: pixelout<=1'b1;
22128: pixelout<=1'b1;
22129: pixelout<=1'b1;
22130: pixelout<=1'b1;
22131: pixelout<=1'b1;
22132: pixelout<=1'b1;
22133: pixelout<=1'b1;
22134: pixelout<=1'b1;
22135: pixelout<=1'b1;
22136: pixelout<=1'b1;
22137: pixelout<=1'b1;
22138: pixelout<=1'b1;
22139: pixelout<=1'b1;
22140: pixelout<=1'b1;
22141: pixelout<=1'b1;
22142: pixelout<=1'b1;
22143: pixelout<=1'b1;
22144: pixelout<=1'b1;
22145: pixelout<=1'b1;
22146: pixelout<=1'b1;
22147: pixelout<=1'b1;
22148: pixelout<=1'b1;
22149: pixelout<=1'b1;
22150: pixelout<=1'b1;
22151: pixelout<=1'b1;
22152: pixelout<=1'b1;
22153: pixelout<=1'b1;
22154: pixelout<=1'b1;
22155: pixelout<=1'b1;
22156: pixelout<=1'b1;
22157: pixelout<=1'b1;
22158: pixelout<=1'b1;
22159: pixelout<=1'b1;
22160: pixelout<=1'b1;
22161: pixelout<=1'b1;
22162: pixelout<=1'b1;
22163: pixelout<=1'b1;
22164: pixelout<=1'b1;
22165: pixelout<=1'b1;
22166: pixelout<=1'b1;
22167: pixelout<=1'b1;
22168: pixelout<=1'b1;
22169: pixelout<=1'b1;
22170: pixelout<=1'b1;
22171: pixelout<=1'b1;
22172: pixelout<=1'b1;
22173: pixelout<=1'b1;
22174: pixelout<=1'b1;
22175: pixelout<=1'b1;
22176: pixelout<=1'b1;
22177: pixelout<=1'b1;
22178: pixelout<=1'b1;
22179: pixelout<=1'b1;
22180: pixelout<=1'b1;
22181: pixelout<=1'b1;
22182: pixelout<=1'b1;
22183: pixelout<=1'b1;
22184: pixelout<=1'b1;
22185: pixelout<=1'b1;
22186: pixelout<=1'b1;
22187: pixelout<=1'b1;
22188: pixelout<=1'b1;
22189: pixelout<=1'b1;
22190: pixelout<=1'b1;
22191: pixelout<=1'b1;
22192: pixelout<=1'b1;
22193: pixelout<=1'b1;
22194: pixelout<=1'b1;
22195: pixelout<=1'b1;
22196: pixelout<=1'b1;
22197: pixelout<=1'b1;
22198: pixelout<=1'b1;
22199: pixelout<=1'b1;
22200: pixelout<=1'b1;
22201: pixelout<=1'b1;
22202: pixelout<=1'b1;
22203: pixelout<=1'b1;
22204: pixelout<=1'b1;
22205: pixelout<=1'b1;
22206: pixelout<=1'b0;
22207: pixelout<=1'b1;
22208: pixelout<=1'b0;
22209: pixelout<=1'b1;
22210: pixelout<=1'b1;
22211: pixelout<=1'b1;
22212: pixelout<=1'b1;
22213: pixelout<=1'b1;
22214: pixelout<=1'b1;
22215: pixelout<=1'b1;
22216: pixelout<=1'b1;
22217: pixelout<=1'b1;
22218: pixelout<=1'b1;
22219: pixelout<=1'b1;
22220: pixelout<=1'b1;
22221: pixelout<=1'b0;
22222: pixelout<=1'b1;
22223: pixelout<=1'b1;
22224: pixelout<=1'b1;
22225: pixelout<=1'b1;
22226: pixelout<=1'b1;
22227: pixelout<=1'b1;
22228: pixelout<=1'b1;
22229: pixelout<=1'b1;
22230: pixelout<=1'b1;
22231: pixelout<=1'b1;
22232: pixelout<=1'b1;
22233: pixelout<=1'b1;
22234: pixelout<=1'b1;
22235: pixelout<=1'b1;
22236: pixelout<=1'b1;
22237: pixelout<=1'b1;
22238: pixelout<=1'b1;
22239: pixelout<=1'b1;
22240: pixelout<=1'b1;
22241: pixelout<=1'b1;
22242: pixelout<=1'b1;
22243: pixelout<=1'b1;
22244: pixelout<=1'b1;
22245: pixelout<=1'b1;
22246: pixelout<=1'b1;
22247: pixelout<=1'b1;
22248: pixelout<=1'b1;
22249: pixelout<=1'b1;
22250: pixelout<=1'b1;
22251: pixelout<=1'b1;
22252: pixelout<=1'b1;
22253: pixelout<=1'b1;
22254: pixelout<=1'b1;
22255: pixelout<=1'b1;
22256: pixelout<=1'b1;
22257: pixelout<=1'b1;
22258: pixelout<=1'b1;
22259: pixelout<=1'b1;
22260: pixelout<=1'b1;
22261: pixelout<=1'b1;
22262: pixelout<=1'b1;
22263: pixelout<=1'b1;
22264: pixelout<=1'b1;
22265: pixelout<=1'b1;
22266: pixelout<=1'b1;
22267: pixelout<=1'b1;
22268: pixelout<=1'b1;
22269: pixelout<=1'b1;
22270: pixelout<=1'b1;
22271: pixelout<=1'b1;
22272: pixelout<=1'b1;
22273: pixelout<=1'b1;
22274: pixelout<=1'b1;
22275: pixelout<=1'b1;
22276: pixelout<=1'b1;
22277: pixelout<=1'b1;
22278: pixelout<=1'b1;
22279: pixelout<=1'b1;
22280: pixelout<=1'b1;
22281: pixelout<=1'b1;
22282: pixelout<=1'b1;
22283: pixelout<=1'b1;
22284: pixelout<=1'b1;
22285: pixelout<=1'b1;
22286: pixelout<=1'b1;
22287: pixelout<=1'b1;
22288: pixelout<=1'b1;
22289: pixelout<=1'b1;
22290: pixelout<=1'b1;
22291: pixelout<=1'b1;
22292: pixelout<=1'b1;
22293: pixelout<=1'b1;
22294: pixelout<=1'b1;
22295: pixelout<=1'b1;
22296: pixelout<=1'b1;
22297: pixelout<=1'b1;
22298: pixelout<=1'b1;
22299: pixelout<=1'b1;
22300: pixelout<=1'b1;
22301: pixelout<=1'b1;
22302: pixelout<=1'b1;
22303: pixelout<=1'b1;
22304: pixelout<=1'b1;
22305: pixelout<=1'b1;
22306: pixelout<=1'b1;
22307: pixelout<=1'b1;
22308: pixelout<=1'b1;
22309: pixelout<=1'b1;
22310: pixelout<=1'b1;
22311: pixelout<=1'b1;
22312: pixelout<=1'b1;
22313: pixelout<=1'b1;
22314: pixelout<=1'b1;
22315: pixelout<=1'b1;
22316: pixelout<=1'b1;
22317: pixelout<=1'b1;
22318: pixelout<=1'b1;
22319: pixelout<=1'b1;
22320: pixelout<=1'b1;
22321: pixelout<=1'b1;
22322: pixelout<=1'b1;
22323: pixelout<=1'b1;
22324: pixelout<=1'b1;
22325: pixelout<=1'b1;
22326: pixelout<=1'b1;
22327: pixelout<=1'b1;
22328: pixelout<=1'b1;
22329: pixelout<=1'b1;
22330: pixelout<=1'b1;
22331: pixelout<=1'b1;
22332: pixelout<=1'b1;
22333: pixelout<=1'b1;
22334: pixelout<=1'b1;
22335: pixelout<=1'b1;
22336: pixelout<=1'b1;
22337: pixelout<=1'b1;
22338: pixelout<=1'b1;
22339: pixelout<=1'b1;
22340: pixelout<=1'b1;
22341: pixelout<=1'b1;
22342: pixelout<=1'b1;
22343: pixelout<=1'b1;
22344: pixelout<=1'b1;
22345: pixelout<=1'b1;
22346: pixelout<=1'b1;
22347: pixelout<=1'b1;
22348: pixelout<=1'b1;
22349: pixelout<=1'b1;
22350: pixelout<=1'b1;
22351: pixelout<=1'b1;
22352: pixelout<=1'b1;
22353: pixelout<=1'b1;
22354: pixelout<=1'b1;
22355: pixelout<=1'b1;
22356: pixelout<=1'b1;
22357: pixelout<=1'b1;
22358: pixelout<=1'b1;
22359: pixelout<=1'b1;
22360: pixelout<=1'b1;
22361: pixelout<=1'b1;
22362: pixelout<=1'b1;
22363: pixelout<=1'b1;
22364: pixelout<=1'b1;
22365: pixelout<=1'b1;
22366: pixelout<=1'b1;
22367: pixelout<=1'b1;
22368: pixelout<=1'b1;
22369: pixelout<=1'b1;
22370: pixelout<=1'b1;
22371: pixelout<=1'b1;
22372: pixelout<=1'b1;
22373: pixelout<=1'b1;
22374: pixelout<=1'b1;
22375: pixelout<=1'b1;
22376: pixelout<=1'b1;
22377: pixelout<=1'b1;
22378: pixelout<=1'b1;
22379: pixelout<=1'b1;
22380: pixelout<=1'b1;
22381: pixelout<=1'b1;
22382: pixelout<=1'b1;
22383: pixelout<=1'b1;
22384: pixelout<=1'b1;
22385: pixelout<=1'b1;
22386: pixelout<=1'b1;
22387: pixelout<=1'b1;
22388: pixelout<=1'b1;
22389: pixelout<=1'b1;
22390: pixelout<=1'b1;
22391: pixelout<=1'b1;
22392: pixelout<=1'b1;
22393: pixelout<=1'b1;
22394: pixelout<=1'b1;
22395: pixelout<=1'b1;
22396: pixelout<=1'b1;
22397: pixelout<=1'b1;
22398: pixelout<=1'b1;
22399: pixelout<=1'b1;
22400: pixelout<=1'b1;
22401: pixelout<=1'b1;
22402: pixelout<=1'b1;
22403: pixelout<=1'b1;
22404: pixelout<=1'b1;
22405: pixelout<=1'b1;
22406: pixelout<=1'b1;
22407: pixelout<=1'b1;
22408: pixelout<=1'b1;
22409: pixelout<=1'b1;
22410: pixelout<=1'b1;
22411: pixelout<=1'b1;
22412: pixelout<=1'b1;
22413: pixelout<=1'b1;
22414: pixelout<=1'b1;
22415: pixelout<=1'b1;
22416: pixelout<=1'b1;
22417: pixelout<=1'b1;
22418: pixelout<=1'b1;
22419: pixelout<=1'b1;
22420: pixelout<=1'b1;
22421: pixelout<=1'b1;
22422: pixelout<=1'b1;
22423: pixelout<=1'b1;
22424: pixelout<=1'b1;
22425: pixelout<=1'b1;
22426: pixelout<=1'b1;
22427: pixelout<=1'b1;
22428: pixelout<=1'b1;
22429: pixelout<=1'b1;
22430: pixelout<=1'b1;
22431: pixelout<=1'b1;
22432: pixelout<=1'b1;
22433: pixelout<=1'b1;
22434: pixelout<=1'b1;
22435: pixelout<=1'b1;
22436: pixelout<=1'b1;
22437: pixelout<=1'b1;
22438: pixelout<=1'b1;
22439: pixelout<=1'b1;
22440: pixelout<=1'b1;
22441: pixelout<=1'b1;
22442: pixelout<=1'b1;
22443: pixelout<=1'b1;
22444: pixelout<=1'b1;
22445: pixelout<=1'b1;
22446: pixelout<=1'b1;
22447: pixelout<=1'b1;
22448: pixelout<=1'b1;
22449: pixelout<=1'b1;
22450: pixelout<=1'b1;
22451: pixelout<=1'b1;
22452: pixelout<=1'b1;
22453: pixelout<=1'b1;
22454: pixelout<=1'b1;
22455: pixelout<=1'b1;
22456: pixelout<=1'b1;
22457: pixelout<=1'b1;
22458: pixelout<=1'b1;
22459: pixelout<=1'b1;
22460: pixelout<=1'b1;
22461: pixelout<=1'b0;
22462: pixelout<=1'b1;
22463: pixelout<=1'b1;
22464: pixelout<=1'b1;
22465: pixelout<=1'b1;
22466: pixelout<=1'b1;
22467: pixelout<=1'b1;
22468: pixelout<=1'b1;
22469: pixelout<=1'b1;
22470: pixelout<=1'b1;
22471: pixelout<=1'b1;
22472: pixelout<=1'b1;
22473: pixelout<=1'b1;
22474: pixelout<=1'b1;
22475: pixelout<=1'b1;
22476: pixelout<=1'b1;
22477: pixelout<=1'b1;
22478: pixelout<=1'b1;
22479: pixelout<=1'b1;
22480: pixelout<=1'b1;
22481: pixelout<=1'b1;
22482: pixelout<=1'b1;
22483: pixelout<=1'b1;
22484: pixelout<=1'b1;
22485: pixelout<=1'b1;
22486: pixelout<=1'b1;
22487: pixelout<=1'b1;
22488: pixelout<=1'b1;
22489: pixelout<=1'b1;
22490: pixelout<=1'b1;
22491: pixelout<=1'b1;
22492: pixelout<=1'b1;
22493: pixelout<=1'b1;
22494: pixelout<=1'b1;
22495: pixelout<=1'b1;
22496: pixelout<=1'b1;
22497: pixelout<=1'b1;
22498: pixelout<=1'b1;
22499: pixelout<=1'b1;
22500: pixelout<=1'b1;
22501: pixelout<=1'b1;
22502: pixelout<=1'b1;
22503: pixelout<=1'b1;
22504: pixelout<=1'b1;
22505: pixelout<=1'b1;
22506: pixelout<=1'b1;
22507: pixelout<=1'b1;
22508: pixelout<=1'b1;
22509: pixelout<=1'b1;
22510: pixelout<=1'b1;
22511: pixelout<=1'b1;
22512: pixelout<=1'b1;
22513: pixelout<=1'b1;
22514: pixelout<=1'b1;
22515: pixelout<=1'b1;
22516: pixelout<=1'b1;
22517: pixelout<=1'b1;
22518: pixelout<=1'b1;
22519: pixelout<=1'b1;
22520: pixelout<=1'b1;
22521: pixelout<=1'b1;
22522: pixelout<=1'b1;
22523: pixelout<=1'b1;
22524: pixelout<=1'b1;
22525: pixelout<=1'b1;
22526: pixelout<=1'b1;
22527: pixelout<=1'b1;
22528: pixelout<=1'b1;
22529: pixelout<=1'b1;
22530: pixelout<=1'b1;
22531: pixelout<=1'b1;
22532: pixelout<=1'b1;
22533: pixelout<=1'b1;
22534: pixelout<=1'b1;
22535: pixelout<=1'b1;
22536: pixelout<=1'b1;
22537: pixelout<=1'b1;
22538: pixelout<=1'b1;
22539: pixelout<=1'b1;
22540: pixelout<=1'b1;
22541: pixelout<=1'b1;
22542: pixelout<=1'b1;
22543: pixelout<=1'b1;
22544: pixelout<=1'b1;
22545: pixelout<=1'b1;
22546: pixelout<=1'b1;
22547: pixelout<=1'b1;
22548: pixelout<=1'b1;
22549: pixelout<=1'b1;
22550: pixelout<=1'b1;
22551: pixelout<=1'b1;
22552: pixelout<=1'b1;
22553: pixelout<=1'b1;
22554: pixelout<=1'b1;
22555: pixelout<=1'b1;
22556: pixelout<=1'b1;
22557: pixelout<=1'b1;
22558: pixelout<=1'b1;
22559: pixelout<=1'b1;
22560: pixelout<=1'b1;
22561: pixelout<=1'b1;
22562: pixelout<=1'b1;
22563: pixelout<=1'b1;
22564: pixelout<=1'b1;
22565: pixelout<=1'b1;
22566: pixelout<=1'b1;
22567: pixelout<=1'b1;
22568: pixelout<=1'b1;
22569: pixelout<=1'b1;
22570: pixelout<=1'b1;
22571: pixelout<=1'b1;
22572: pixelout<=1'b1;
22573: pixelout<=1'b1;
22574: pixelout<=1'b1;
22575: pixelout<=1'b1;
22576: pixelout<=1'b1;
22577: pixelout<=1'b1;
22578: pixelout<=1'b1;
22579: pixelout<=1'b1;
22580: pixelout<=1'b1;
22581: pixelout<=1'b1;
22582: pixelout<=1'b1;
22583: pixelout<=1'b1;
22584: pixelout<=1'b1;
22585: pixelout<=1'b1;
22586: pixelout<=1'b1;
22587: pixelout<=1'b1;
22588: pixelout<=1'b1;
22589: pixelout<=1'b1;
22590: pixelout<=1'b1;
22591: pixelout<=1'b1;
22592: pixelout<=1'b1;
22593: pixelout<=1'b1;
22594: pixelout<=1'b1;
22595: pixelout<=1'b1;
22596: pixelout<=1'b1;
22597: pixelout<=1'b1;
22598: pixelout<=1'b1;
22599: pixelout<=1'b1;
22600: pixelout<=1'b1;
22601: pixelout<=1'b1;
22602: pixelout<=1'b1;
22603: pixelout<=1'b1;
22604: pixelout<=1'b1;
22605: pixelout<=1'b1;
22606: pixelout<=1'b1;
22607: pixelout<=1'b1;
22608: pixelout<=1'b1;
22609: pixelout<=1'b1;
22610: pixelout<=1'b1;
22611: pixelout<=1'b1;
22612: pixelout<=1'b1;
22613: pixelout<=1'b1;
22614: pixelout<=1'b1;
22615: pixelout<=1'b1;
22616: pixelout<=1'b1;
22617: pixelout<=1'b1;
22618: pixelout<=1'b1;
22619: pixelout<=1'b1;
22620: pixelout<=1'b1;
22621: pixelout<=1'b1;
22622: pixelout<=1'b1;
22623: pixelout<=1'b1;
22624: pixelout<=1'b1;
22625: pixelout<=1'b1;
22626: pixelout<=1'b1;
22627: pixelout<=1'b1;
22628: pixelout<=1'b1;
22629: pixelout<=1'b1;
22630: pixelout<=1'b1;
22631: pixelout<=1'b1;
22632: pixelout<=1'b1;
22633: pixelout<=1'b1;
22634: pixelout<=1'b1;
22635: pixelout<=1'b1;
22636: pixelout<=1'b1;
22637: pixelout<=1'b1;
22638: pixelout<=1'b1;
22639: pixelout<=1'b1;
22640: pixelout<=1'b1;
22641: pixelout<=1'b1;
22642: pixelout<=1'b1;
22643: pixelout<=1'b1;
22644: pixelout<=1'b1;
22645: pixelout<=1'b1;
22646: pixelout<=1'b1;
22647: pixelout<=1'b1;
22648: pixelout<=1'b1;
22649: pixelout<=1'b1;
22650: pixelout<=1'b1;
22651: pixelout<=1'b1;
22652: pixelout<=1'b1;
22653: pixelout<=1'b1;
22654: pixelout<=1'b1;
22655: pixelout<=1'b1;
22656: pixelout<=1'b1;
22657: pixelout<=1'b1;
22658: pixelout<=1'b1;
22659: pixelout<=1'b0;
22660: pixelout<=1'b1;
22661: pixelout<=1'b1;
22662: pixelout<=1'b0;
22663: pixelout<=1'b1;
22664: pixelout<=1'b1;
22665: pixelout<=1'b0;
22666: pixelout<=1'b0;
22667: pixelout<=1'b0;
22668: pixelout<=1'b0;
22669: pixelout<=1'b1;
22670: pixelout<=1'b1;
22671: pixelout<=1'b1;
22672: pixelout<=1'b1;
22673: pixelout<=1'b1;
22674: pixelout<=1'b1;
22675: pixelout<=1'b0;
22676: pixelout<=1'b0;
22677: pixelout<=1'b1;
22678: pixelout<=1'b1;
22679: pixelout<=1'b1;
22680: pixelout<=1'b1;
22681: pixelout<=1'b1;
22682: pixelout<=1'b1;
22683: pixelout<=1'b1;
22684: pixelout<=1'b0;
22685: pixelout<=1'b0;
22686: pixelout<=1'b1;
22687: pixelout<=1'b1;
22688: pixelout<=1'b1;
22689: pixelout<=1'b1;
22690: pixelout<=1'b0;
22691: pixelout<=1'b0;
22692: pixelout<=1'b1;
22693: pixelout<=1'b1;
22694: pixelout<=1'b1;
22695: pixelout<=1'b0;
22696: pixelout<=1'b0;
22697: pixelout<=1'b0;
22698: pixelout<=1'b1;
22699: pixelout<=1'b1;
22700: pixelout<=1'b1;
22701: pixelout<=1'b0;
22702: pixelout<=1'b1;
22703: pixelout<=1'b1;
22704: pixelout<=1'b1;
22705: pixelout<=1'b1;
22706: pixelout<=1'b1;
22707: pixelout<=1'b1;
22708: pixelout<=1'b1;
22709: pixelout<=1'b1;
22710: pixelout<=1'b1;
22711: pixelout<=1'b1;
22712: pixelout<=1'b1;
22713: pixelout<=1'b1;
22714: pixelout<=1'b1;
22715: pixelout<=1'b1;
22716: pixelout<=1'b1;
22717: pixelout<=1'b1;
22718: pixelout<=1'b1;
22719: pixelout<=1'b1;
22720: pixelout<=1'b1;
22721: pixelout<=1'b1;
22722: pixelout<=1'b1;
22723: pixelout<=1'b1;
22724: pixelout<=1'b1;
22725: pixelout<=1'b1;
22726: pixelout<=1'b1;
22727: pixelout<=1'b1;
22728: pixelout<=1'b1;
22729: pixelout<=1'b1;
22730: pixelout<=1'b1;
22731: pixelout<=1'b1;
22732: pixelout<=1'b1;
22733: pixelout<=1'b1;
22734: pixelout<=1'b1;
22735: pixelout<=1'b1;
22736: pixelout<=1'b1;
22737: pixelout<=1'b1;
22738: pixelout<=1'b1;
22739: pixelout<=1'b1;
22740: pixelout<=1'b1;
22741: pixelout<=1'b1;
22742: pixelout<=1'b1;
22743: pixelout<=1'b1;
22744: pixelout<=1'b1;
22745: pixelout<=1'b1;
22746: pixelout<=1'b1;
22747: pixelout<=1'b1;
22748: pixelout<=1'b1;
22749: pixelout<=1'b1;
22750: pixelout<=1'b1;
22751: pixelout<=1'b1;
22752: pixelout<=1'b1;
22753: pixelout<=1'b1;
22754: pixelout<=1'b1;
22755: pixelout<=1'b1;
22756: pixelout<=1'b1;
22757: pixelout<=1'b1;
22758: pixelout<=1'b1;
22759: pixelout<=1'b1;
22760: pixelout<=1'b1;
22761: pixelout<=1'b1;
22762: pixelout<=1'b1;
22763: pixelout<=1'b1;
22764: pixelout<=1'b1;
22765: pixelout<=1'b1;
22766: pixelout<=1'b1;
22767: pixelout<=1'b1;
22768: pixelout<=1'b1;
22769: pixelout<=1'b1;
22770: pixelout<=1'b1;
22771: pixelout<=1'b1;
22772: pixelout<=1'b1;
22773: pixelout<=1'b1;
22774: pixelout<=1'b1;
22775: pixelout<=1'b1;
22776: pixelout<=1'b1;
22777: pixelout<=1'b1;
22778: pixelout<=1'b1;
22779: pixelout<=1'b1;
22780: pixelout<=1'b1;
22781: pixelout<=1'b1;
22782: pixelout<=1'b1;
22783: pixelout<=1'b1;
22784: pixelout<=1'b1;
22785: pixelout<=1'b1;
22786: pixelout<=1'b1;
22787: pixelout<=1'b1;
22788: pixelout<=1'b1;
22789: pixelout<=1'b1;
22790: pixelout<=1'b1;
22791: pixelout<=1'b1;
22792: pixelout<=1'b1;
22793: pixelout<=1'b1;
22794: pixelout<=1'b1;
22795: pixelout<=1'b1;
22796: pixelout<=1'b1;
22797: pixelout<=1'b1;
22798: pixelout<=1'b1;
22799: pixelout<=1'b1;
22800: pixelout<=1'b1;
22801: pixelout<=1'b1;
22802: pixelout<=1'b1;
22803: pixelout<=1'b1;
22804: pixelout<=1'b1;
22805: pixelout<=1'b1;
22806: pixelout<=1'b1;
22807: pixelout<=1'b1;
22808: pixelout<=1'b1;
22809: pixelout<=1'b1;
22810: pixelout<=1'b1;
22811: pixelout<=1'b1;
22812: pixelout<=1'b1;
22813: pixelout<=1'b1;
22814: pixelout<=1'b1;
22815: pixelout<=1'b1;
22816: pixelout<=1'b1;
22817: pixelout<=1'b1;
22818: pixelout<=1'b1;
22819: pixelout<=1'b1;
22820: pixelout<=1'b1;
22821: pixelout<=1'b1;
22822: pixelout<=1'b1;
22823: pixelout<=1'b1;
22824: pixelout<=1'b1;
22825: pixelout<=1'b1;
22826: pixelout<=1'b1;
22827: pixelout<=1'b1;
22828: pixelout<=1'b1;
22829: pixelout<=1'b1;
22830: pixelout<=1'b1;
22831: pixelout<=1'b1;
22832: pixelout<=1'b1;
22833: pixelout<=1'b1;
22834: pixelout<=1'b1;
22835: pixelout<=1'b1;
22836: pixelout<=1'b1;
22837: pixelout<=1'b1;
22838: pixelout<=1'b1;
22839: pixelout<=1'b1;
22840: pixelout<=1'b1;
22841: pixelout<=1'b1;
22842: pixelout<=1'b1;
22843: pixelout<=1'b1;
22844: pixelout<=1'b1;
22845: pixelout<=1'b1;
22846: pixelout<=1'b1;
22847: pixelout<=1'b1;
22848: pixelout<=1'b1;
22849: pixelout<=1'b1;
22850: pixelout<=1'b1;
22851: pixelout<=1'b1;
22852: pixelout<=1'b1;
22853: pixelout<=1'b1;
22854: pixelout<=1'b1;
22855: pixelout<=1'b1;
22856: pixelout<=1'b1;
22857: pixelout<=1'b1;
22858: pixelout<=1'b1;
22859: pixelout<=1'b1;
22860: pixelout<=1'b1;
22861: pixelout<=1'b1;
22862: pixelout<=1'b1;
22863: pixelout<=1'b1;
22864: pixelout<=1'b1;
22865: pixelout<=1'b1;
22866: pixelout<=1'b1;
22867: pixelout<=1'b1;
22868: pixelout<=1'b1;
22869: pixelout<=1'b1;
22870: pixelout<=1'b1;
22871: pixelout<=1'b1;
22872: pixelout<=1'b1;
22873: pixelout<=1'b1;
22874: pixelout<=1'b1;
22875: pixelout<=1'b1;
22876: pixelout<=1'b1;
22877: pixelout<=1'b1;
22878: pixelout<=1'b1;
22879: pixelout<=1'b1;
22880: pixelout<=1'b1;
22881: pixelout<=1'b1;
22882: pixelout<=1'b1;
22883: pixelout<=1'b1;
22884: pixelout<=1'b1;
22885: pixelout<=1'b1;
22886: pixelout<=1'b1;
22887: pixelout<=1'b1;
22888: pixelout<=1'b1;
22889: pixelout<=1'b1;
22890: pixelout<=1'b1;
22891: pixelout<=1'b1;
22892: pixelout<=1'b1;
22893: pixelout<=1'b1;
22894: pixelout<=1'b1;
22895: pixelout<=1'b1;
22896: pixelout<=1'b1;
22897: pixelout<=1'b1;
22898: pixelout<=1'b1;
22899: pixelout<=1'b0;
22900: pixelout<=1'b1;
22901: pixelout<=1'b1;
22902: pixelout<=1'b0;
22903: pixelout<=1'b1;
22904: pixelout<=1'b1;
22905: pixelout<=1'b0;
22906: pixelout<=1'b1;
22907: pixelout<=1'b1;
22908: pixelout<=1'b1;
22909: pixelout<=1'b1;
22910: pixelout<=1'b1;
22911: pixelout<=1'b1;
22912: pixelout<=1'b1;
22913: pixelout<=1'b1;
22914: pixelout<=1'b1;
22915: pixelout<=1'b1;
22916: pixelout<=1'b1;
22917: pixelout<=1'b1;
22918: pixelout<=1'b0;
22919: pixelout<=1'b1;
22920: pixelout<=1'b1;
22921: pixelout<=1'b1;
22922: pixelout<=1'b1;
22923: pixelout<=1'b1;
22924: pixelout<=1'b1;
22925: pixelout<=1'b1;
22926: pixelout<=1'b0;
22927: pixelout<=1'b1;
22928: pixelout<=1'b0;
22929: pixelout<=1'b1;
22930: pixelout<=1'b1;
22931: pixelout<=1'b1;
22932: pixelout<=1'b1;
22933: pixelout<=1'b1;
22934: pixelout<=1'b1;
22935: pixelout<=1'b1;
22936: pixelout<=1'b1;
22937: pixelout<=1'b1;
22938: pixelout<=1'b1;
22939: pixelout<=1'b0;
22940: pixelout<=1'b1;
22941: pixelout<=1'b0;
22942: pixelout<=1'b1;
22943: pixelout<=1'b1;
22944: pixelout<=1'b1;
22945: pixelout<=1'b1;
22946: pixelout<=1'b1;
22947: pixelout<=1'b1;
22948: pixelout<=1'b1;
22949: pixelout<=1'b1;
22950: pixelout<=1'b1;
22951: pixelout<=1'b1;
22952: pixelout<=1'b1;
22953: pixelout<=1'b1;
22954: pixelout<=1'b1;
22955: pixelout<=1'b1;
22956: pixelout<=1'b1;
22957: pixelout<=1'b1;
22958: pixelout<=1'b1;
22959: pixelout<=1'b1;
22960: pixelout<=1'b1;
22961: pixelout<=1'b1;
22962: pixelout<=1'b1;
22963: pixelout<=1'b1;
22964: pixelout<=1'b1;
22965: pixelout<=1'b1;
22966: pixelout<=1'b1;
22967: pixelout<=1'b1;
22968: pixelout<=1'b1;
22969: pixelout<=1'b1;
22970: pixelout<=1'b1;
22971: pixelout<=1'b1;
22972: pixelout<=1'b1;
22973: pixelout<=1'b1;
22974: pixelout<=1'b1;
22975: pixelout<=1'b1;
22976: pixelout<=1'b1;
22977: pixelout<=1'b1;
22978: pixelout<=1'b1;
22979: pixelout<=1'b1;
22980: pixelout<=1'b1;
22981: pixelout<=1'b1;
22982: pixelout<=1'b1;
22983: pixelout<=1'b1;
22984: pixelout<=1'b1;
22985: pixelout<=1'b1;
22986: pixelout<=1'b1;
22987: pixelout<=1'b1;
22988: pixelout<=1'b1;
22989: pixelout<=1'b1;
22990: pixelout<=1'b1;
22991: pixelout<=1'b1;
22992: pixelout<=1'b1;
22993: pixelout<=1'b1;
22994: pixelout<=1'b1;
22995: pixelout<=1'b1;
22996: pixelout<=1'b1;
22997: pixelout<=1'b1;
22998: pixelout<=1'b1;
22999: pixelout<=1'b1;
23000: pixelout<=1'b1;
23001: pixelout<=1'b1;
23002: pixelout<=1'b1;
23003: pixelout<=1'b1;
23004: pixelout<=1'b1;
23005: pixelout<=1'b1;
23006: pixelout<=1'b1;
23007: pixelout<=1'b1;
23008: pixelout<=1'b1;
23009: pixelout<=1'b1;
23010: pixelout<=1'b1;
23011: pixelout<=1'b1;
23012: pixelout<=1'b1;
23013: pixelout<=1'b1;
23014: pixelout<=1'b1;
23015: pixelout<=1'b1;
23016: pixelout<=1'b1;
23017: pixelout<=1'b1;
23018: pixelout<=1'b1;
23019: pixelout<=1'b1;
23020: pixelout<=1'b1;
23021: pixelout<=1'b1;
23022: pixelout<=1'b1;
23023: pixelout<=1'b1;
23024: pixelout<=1'b1;
23025: pixelout<=1'b1;
23026: pixelout<=1'b1;
23027: pixelout<=1'b1;
23028: pixelout<=1'b1;
23029: pixelout<=1'b1;
23030: pixelout<=1'b1;
23031: pixelout<=1'b1;
23032: pixelout<=1'b1;
23033: pixelout<=1'b1;
23034: pixelout<=1'b1;
23035: pixelout<=1'b1;
23036: pixelout<=1'b1;
23037: pixelout<=1'b1;
23038: pixelout<=1'b1;
23039: pixelout<=1'b1;
23040: pixelout<=1'b1;
23041: pixelout<=1'b1;
23042: pixelout<=1'b1;
23043: pixelout<=1'b1;
23044: pixelout<=1'b1;
23045: pixelout<=1'b1;
23046: pixelout<=1'b1;
23047: pixelout<=1'b1;
23048: pixelout<=1'b1;
23049: pixelout<=1'b1;
23050: pixelout<=1'b1;
23051: pixelout<=1'b1;
23052: pixelout<=1'b1;
23053: pixelout<=1'b1;
23054: pixelout<=1'b1;
23055: pixelout<=1'b1;
23056: pixelout<=1'b1;
23057: pixelout<=1'b1;
23058: pixelout<=1'b1;
23059: pixelout<=1'b1;
23060: pixelout<=1'b1;
23061: pixelout<=1'b1;
23062: pixelout<=1'b1;
23063: pixelout<=1'b1;
23064: pixelout<=1'b1;
23065: pixelout<=1'b1;
23066: pixelout<=1'b1;
23067: pixelout<=1'b1;
23068: pixelout<=1'b1;
23069: pixelout<=1'b1;
23070: pixelout<=1'b1;
23071: pixelout<=1'b1;
23072: pixelout<=1'b1;
23073: pixelout<=1'b1;
23074: pixelout<=1'b1;
23075: pixelout<=1'b1;
23076: pixelout<=1'b1;
23077: pixelout<=1'b1;
23078: pixelout<=1'b1;
23079: pixelout<=1'b1;
23080: pixelout<=1'b1;
23081: pixelout<=1'b1;
23082: pixelout<=1'b1;
23083: pixelout<=1'b1;
23084: pixelout<=1'b1;
23085: pixelout<=1'b1;
23086: pixelout<=1'b1;
23087: pixelout<=1'b1;
23088: pixelout<=1'b1;
23089: pixelout<=1'b1;
23090: pixelout<=1'b1;
23091: pixelout<=1'b1;
23092: pixelout<=1'b1;
23093: pixelout<=1'b1;
23094: pixelout<=1'b1;
23095: pixelout<=1'b1;
23096: pixelout<=1'b1;
23097: pixelout<=1'b1;
23098: pixelout<=1'b1;
23099: pixelout<=1'b1;
23100: pixelout<=1'b1;
23101: pixelout<=1'b1;
23102: pixelout<=1'b1;
23103: pixelout<=1'b1;
23104: pixelout<=1'b1;
23105: pixelout<=1'b1;
23106: pixelout<=1'b1;
23107: pixelout<=1'b1;
23108: pixelout<=1'b1;
23109: pixelout<=1'b1;
23110: pixelout<=1'b1;
23111: pixelout<=1'b1;
23112: pixelout<=1'b1;
23113: pixelout<=1'b1;
23114: pixelout<=1'b1;
23115: pixelout<=1'b1;
23116: pixelout<=1'b1;
23117: pixelout<=1'b1;
23118: pixelout<=1'b1;
23119: pixelout<=1'b1;
23120: pixelout<=1'b1;
23121: pixelout<=1'b1;
23122: pixelout<=1'b1;
23123: pixelout<=1'b1;
23124: pixelout<=1'b1;
23125: pixelout<=1'b1;
23126: pixelout<=1'b1;
23127: pixelout<=1'b1;
23128: pixelout<=1'b1;
23129: pixelout<=1'b1;
23130: pixelout<=1'b1;
23131: pixelout<=1'b1;
23132: pixelout<=1'b1;
23133: pixelout<=1'b1;
23134: pixelout<=1'b1;
23135: pixelout<=1'b1;
23136: pixelout<=1'b1;
23137: pixelout<=1'b1;
23138: pixelout<=1'b1;
23139: pixelout<=1'b0;
23140: pixelout<=1'b1;
23141: pixelout<=1'b1;
23142: pixelout<=1'b0;
23143: pixelout<=1'b1;
23144: pixelout<=1'b1;
23145: pixelout<=1'b1;
23146: pixelout<=1'b0;
23147: pixelout<=1'b0;
23148: pixelout<=1'b1;
23149: pixelout<=1'b1;
23150: pixelout<=1'b1;
23151: pixelout<=1'b1;
23152: pixelout<=1'b1;
23153: pixelout<=1'b1;
23154: pixelout<=1'b1;
23155: pixelout<=1'b1;
23156: pixelout<=1'b1;
23157: pixelout<=1'b1;
23158: pixelout<=1'b0;
23159: pixelout<=1'b1;
23160: pixelout<=1'b1;
23161: pixelout<=1'b1;
23162: pixelout<=1'b1;
23163: pixelout<=1'b1;
23164: pixelout<=1'b1;
23165: pixelout<=1'b1;
23166: pixelout<=1'b0;
23167: pixelout<=1'b1;
23168: pixelout<=1'b0;
23169: pixelout<=1'b1;
23170: pixelout<=1'b1;
23171: pixelout<=1'b1;
23172: pixelout<=1'b1;
23173: pixelout<=1'b1;
23174: pixelout<=1'b1;
23175: pixelout<=1'b1;
23176: pixelout<=1'b1;
23177: pixelout<=1'b1;
23178: pixelout<=1'b1;
23179: pixelout<=1'b0;
23180: pixelout<=1'b1;
23181: pixelout<=1'b1;
23182: pixelout<=1'b1;
23183: pixelout<=1'b1;
23184: pixelout<=1'b1;
23185: pixelout<=1'b1;
23186: pixelout<=1'b1;
23187: pixelout<=1'b1;
23188: pixelout<=1'b1;
23189: pixelout<=1'b1;
23190: pixelout<=1'b1;
23191: pixelout<=1'b1;
23192: pixelout<=1'b1;
23193: pixelout<=1'b1;
23194: pixelout<=1'b1;
23195: pixelout<=1'b1;
23196: pixelout<=1'b1;
23197: pixelout<=1'b1;
23198: pixelout<=1'b1;
23199: pixelout<=1'b1;
23200: pixelout<=1'b1;
23201: pixelout<=1'b1;
23202: pixelout<=1'b1;
23203: pixelout<=1'b1;
23204: pixelout<=1'b1;
23205: pixelout<=1'b1;
23206: pixelout<=1'b1;
23207: pixelout<=1'b1;
23208: pixelout<=1'b1;
23209: pixelout<=1'b1;
23210: pixelout<=1'b1;
23211: pixelout<=1'b1;
23212: pixelout<=1'b1;
23213: pixelout<=1'b1;
23214: pixelout<=1'b1;
23215: pixelout<=1'b1;
23216: pixelout<=1'b1;
23217: pixelout<=1'b1;
23218: pixelout<=1'b1;
23219: pixelout<=1'b1;
23220: pixelout<=1'b1;
23221: pixelout<=1'b1;
23222: pixelout<=1'b1;
23223: pixelout<=1'b1;
23224: pixelout<=1'b1;
23225: pixelout<=1'b1;
23226: pixelout<=1'b1;
23227: pixelout<=1'b1;
23228: pixelout<=1'b1;
23229: pixelout<=1'b1;
23230: pixelout<=1'b1;
23231: pixelout<=1'b1;
23232: pixelout<=1'b1;
23233: pixelout<=1'b1;
23234: pixelout<=1'b1;
23235: pixelout<=1'b1;
23236: pixelout<=1'b1;
23237: pixelout<=1'b1;
23238: pixelout<=1'b1;
23239: pixelout<=1'b1;
23240: pixelout<=1'b1;
23241: pixelout<=1'b1;
23242: pixelout<=1'b1;
23243: pixelout<=1'b1;
23244: pixelout<=1'b1;
23245: pixelout<=1'b1;
23246: pixelout<=1'b1;
23247: pixelout<=1'b1;
23248: pixelout<=1'b1;
23249: pixelout<=1'b1;
23250: pixelout<=1'b1;
23251: pixelout<=1'b1;
23252: pixelout<=1'b1;
23253: pixelout<=1'b1;
23254: pixelout<=1'b1;
23255: pixelout<=1'b1;
23256: pixelout<=1'b1;
23257: pixelout<=1'b1;
23258: pixelout<=1'b1;
23259: pixelout<=1'b1;
23260: pixelout<=1'b1;
23261: pixelout<=1'b1;
23262: pixelout<=1'b1;
23263: pixelout<=1'b1;
23264: pixelout<=1'b1;
23265: pixelout<=1'b1;
23266: pixelout<=1'b1;
23267: pixelout<=1'b1;
23268: pixelout<=1'b1;
23269: pixelout<=1'b1;
23270: pixelout<=1'b1;
23271: pixelout<=1'b1;
23272: pixelout<=1'b1;
23273: pixelout<=1'b1;
23274: pixelout<=1'b1;
23275: pixelout<=1'b1;
23276: pixelout<=1'b1;
23277: pixelout<=1'b1;
23278: pixelout<=1'b1;
23279: pixelout<=1'b1;
23280: pixelout<=1'b1;
23281: pixelout<=1'b1;
23282: pixelout<=1'b1;
23283: pixelout<=1'b1;
23284: pixelout<=1'b1;
23285: pixelout<=1'b1;
23286: pixelout<=1'b1;
23287: pixelout<=1'b1;
23288: pixelout<=1'b1;
23289: pixelout<=1'b1;
23290: pixelout<=1'b1;
23291: pixelout<=1'b1;
23292: pixelout<=1'b1;
23293: pixelout<=1'b1;
23294: pixelout<=1'b1;
23295: pixelout<=1'b1;
23296: pixelout<=1'b1;
23297: pixelout<=1'b1;
23298: pixelout<=1'b1;
23299: pixelout<=1'b1;
23300: pixelout<=1'b1;
23301: pixelout<=1'b1;
23302: pixelout<=1'b1;
23303: pixelout<=1'b1;
23304: pixelout<=1'b1;
23305: pixelout<=1'b1;
23306: pixelout<=1'b1;
23307: pixelout<=1'b1;
23308: pixelout<=1'b1;
23309: pixelout<=1'b1;
23310: pixelout<=1'b1;
23311: pixelout<=1'b1;
23312: pixelout<=1'b1;
23313: pixelout<=1'b1;
23314: pixelout<=1'b1;
23315: pixelout<=1'b1;
23316: pixelout<=1'b1;
23317: pixelout<=1'b1;
23318: pixelout<=1'b1;
23319: pixelout<=1'b1;
23320: pixelout<=1'b1;
23321: pixelout<=1'b1;
23322: pixelout<=1'b1;
23323: pixelout<=1'b1;
23324: pixelout<=1'b1;
23325: pixelout<=1'b1;
23326: pixelout<=1'b1;
23327: pixelout<=1'b1;
23328: pixelout<=1'b1;
23329: pixelout<=1'b1;
23330: pixelout<=1'b1;
23331: pixelout<=1'b1;
23332: pixelout<=1'b1;
23333: pixelout<=1'b1;
23334: pixelout<=1'b1;
23335: pixelout<=1'b1;
23336: pixelout<=1'b1;
23337: pixelout<=1'b1;
23338: pixelout<=1'b1;
23339: pixelout<=1'b1;
23340: pixelout<=1'b1;
23341: pixelout<=1'b1;
23342: pixelout<=1'b1;
23343: pixelout<=1'b1;
23344: pixelout<=1'b1;
23345: pixelout<=1'b1;
23346: pixelout<=1'b1;
23347: pixelout<=1'b1;
23348: pixelout<=1'b1;
23349: pixelout<=1'b1;
23350: pixelout<=1'b1;
23351: pixelout<=1'b1;
23352: pixelout<=1'b1;
23353: pixelout<=1'b1;
23354: pixelout<=1'b1;
23355: pixelout<=1'b1;
23356: pixelout<=1'b1;
23357: pixelout<=1'b1;
23358: pixelout<=1'b1;
23359: pixelout<=1'b1;
23360: pixelout<=1'b1;
23361: pixelout<=1'b1;
23362: pixelout<=1'b1;
23363: pixelout<=1'b1;
23364: pixelout<=1'b1;
23365: pixelout<=1'b1;
23366: pixelout<=1'b1;
23367: pixelout<=1'b1;
23368: pixelout<=1'b1;
23369: pixelout<=1'b1;
23370: pixelout<=1'b1;
23371: pixelout<=1'b1;
23372: pixelout<=1'b1;
23373: pixelout<=1'b1;
23374: pixelout<=1'b1;
23375: pixelout<=1'b1;
23376: pixelout<=1'b1;
23377: pixelout<=1'b1;
23378: pixelout<=1'b1;
23379: pixelout<=1'b0;
23380: pixelout<=1'b1;
23381: pixelout<=1'b1;
23382: pixelout<=1'b0;
23383: pixelout<=1'b1;
23384: pixelout<=1'b1;
23385: pixelout<=1'b1;
23386: pixelout<=1'b1;
23387: pixelout<=1'b1;
23388: pixelout<=1'b0;
23389: pixelout<=1'b1;
23390: pixelout<=1'b1;
23391: pixelout<=1'b1;
23392: pixelout<=1'b1;
23393: pixelout<=1'b1;
23394: pixelout<=1'b1;
23395: pixelout<=1'b1;
23396: pixelout<=1'b1;
23397: pixelout<=1'b1;
23398: pixelout<=1'b0;
23399: pixelout<=1'b1;
23400: pixelout<=1'b1;
23401: pixelout<=1'b1;
23402: pixelout<=1'b0;
23403: pixelout<=1'b1;
23404: pixelout<=1'b1;
23405: pixelout<=1'b1;
23406: pixelout<=1'b0;
23407: pixelout<=1'b1;
23408: pixelout<=1'b0;
23409: pixelout<=1'b1;
23410: pixelout<=1'b1;
23411: pixelout<=1'b1;
23412: pixelout<=1'b1;
23413: pixelout<=1'b1;
23414: pixelout<=1'b1;
23415: pixelout<=1'b1;
23416: pixelout<=1'b1;
23417: pixelout<=1'b1;
23418: pixelout<=1'b1;
23419: pixelout<=1'b0;
23420: pixelout<=1'b1;
23421: pixelout<=1'b0;
23422: pixelout<=1'b1;
23423: pixelout<=1'b1;
23424: pixelout<=1'b1;
23425: pixelout<=1'b1;
23426: pixelout<=1'b1;
23427: pixelout<=1'b1;
23428: pixelout<=1'b1;
23429: pixelout<=1'b1;
23430: pixelout<=1'b1;
23431: pixelout<=1'b1;
23432: pixelout<=1'b1;
23433: pixelout<=1'b1;
23434: pixelout<=1'b1;
23435: pixelout<=1'b1;
23436: pixelout<=1'b1;
23437: pixelout<=1'b1;
23438: pixelout<=1'b1;
23439: pixelout<=1'b1;
23440: pixelout<=1'b1;
23441: pixelout<=1'b1;
23442: pixelout<=1'b1;
23443: pixelout<=1'b1;
23444: pixelout<=1'b1;
23445: pixelout<=1'b1;
23446: pixelout<=1'b1;
23447: pixelout<=1'b1;
23448: pixelout<=1'b1;
23449: pixelout<=1'b1;
23450: pixelout<=1'b1;
23451: pixelout<=1'b1;
23452: pixelout<=1'b1;
23453: pixelout<=1'b1;
23454: pixelout<=1'b1;
23455: pixelout<=1'b1;
23456: pixelout<=1'b1;
23457: pixelout<=1'b1;
23458: pixelout<=1'b1;
23459: pixelout<=1'b1;
23460: pixelout<=1'b1;
23461: pixelout<=1'b1;
23462: pixelout<=1'b1;
23463: pixelout<=1'b1;
23464: pixelout<=1'b1;
23465: pixelout<=1'b1;
23466: pixelout<=1'b1;
23467: pixelout<=1'b1;
23468: pixelout<=1'b1;
23469: pixelout<=1'b1;
23470: pixelout<=1'b1;
23471: pixelout<=1'b1;
23472: pixelout<=1'b1;
23473: pixelout<=1'b1;
23474: pixelout<=1'b1;
23475: pixelout<=1'b1;
23476: pixelout<=1'b1;
23477: pixelout<=1'b1;
23478: pixelout<=1'b1;
23479: pixelout<=1'b1;
23480: pixelout<=1'b1;
23481: pixelout<=1'b1;
23482: pixelout<=1'b1;
23483: pixelout<=1'b1;
23484: pixelout<=1'b1;
23485: pixelout<=1'b1;
23486: pixelout<=1'b1;
23487: pixelout<=1'b1;
23488: pixelout<=1'b1;
23489: pixelout<=1'b1;
23490: pixelout<=1'b1;
23491: pixelout<=1'b1;
23492: pixelout<=1'b1;
23493: pixelout<=1'b1;
23494: pixelout<=1'b1;
23495: pixelout<=1'b1;
23496: pixelout<=1'b1;
23497: pixelout<=1'b1;
23498: pixelout<=1'b1;
23499: pixelout<=1'b1;
23500: pixelout<=1'b1;
23501: pixelout<=1'b1;
23502: pixelout<=1'b1;
23503: pixelout<=1'b1;
23504: pixelout<=1'b1;
23505: pixelout<=1'b1;
23506: pixelout<=1'b1;
23507: pixelout<=1'b1;
23508: pixelout<=1'b1;
23509: pixelout<=1'b1;
23510: pixelout<=1'b1;
23511: pixelout<=1'b1;
23512: pixelout<=1'b1;
23513: pixelout<=1'b1;
23514: pixelout<=1'b1;
23515: pixelout<=1'b1;
23516: pixelout<=1'b1;
23517: pixelout<=1'b1;
23518: pixelout<=1'b1;
23519: pixelout<=1'b1;
23520: pixelout<=1'b1;
23521: pixelout<=1'b1;
23522: pixelout<=1'b1;
23523: pixelout<=1'b1;
23524: pixelout<=1'b1;
23525: pixelout<=1'b1;
23526: pixelout<=1'b1;
23527: pixelout<=1'b1;
23528: pixelout<=1'b1;
23529: pixelout<=1'b1;
23530: pixelout<=1'b1;
23531: pixelout<=1'b1;
23532: pixelout<=1'b1;
23533: pixelout<=1'b1;
23534: pixelout<=1'b1;
23535: pixelout<=1'b1;
23536: pixelout<=1'b1;
23537: pixelout<=1'b1;
23538: pixelout<=1'b1;
23539: pixelout<=1'b1;
23540: pixelout<=1'b1;
23541: pixelout<=1'b1;
23542: pixelout<=1'b1;
23543: pixelout<=1'b1;
23544: pixelout<=1'b1;
23545: pixelout<=1'b1;
23546: pixelout<=1'b1;
23547: pixelout<=1'b1;
23548: pixelout<=1'b1;
23549: pixelout<=1'b1;
23550: pixelout<=1'b1;
23551: pixelout<=1'b1;
23552: pixelout<=1'b1;
23553: pixelout<=1'b1;
23554: pixelout<=1'b1;
23555: pixelout<=1'b1;
23556: pixelout<=1'b1;
23557: pixelout<=1'b1;
23558: pixelout<=1'b1;
23559: pixelout<=1'b1;
23560: pixelout<=1'b1;
23561: pixelout<=1'b1;
23562: pixelout<=1'b1;
23563: pixelout<=1'b1;
23564: pixelout<=1'b1;
23565: pixelout<=1'b1;
23566: pixelout<=1'b1;
23567: pixelout<=1'b1;
23568: pixelout<=1'b1;
23569: pixelout<=1'b1;
23570: pixelout<=1'b1;
23571: pixelout<=1'b1;
23572: pixelout<=1'b1;
23573: pixelout<=1'b1;
23574: pixelout<=1'b1;
23575: pixelout<=1'b1;
23576: pixelout<=1'b1;
23577: pixelout<=1'b1;
23578: pixelout<=1'b1;
23579: pixelout<=1'b1;
23580: pixelout<=1'b1;
23581: pixelout<=1'b1;
23582: pixelout<=1'b1;
23583: pixelout<=1'b1;
23584: pixelout<=1'b1;
23585: pixelout<=1'b1;
23586: pixelout<=1'b1;
23587: pixelout<=1'b1;
23588: pixelout<=1'b1;
23589: pixelout<=1'b1;
23590: pixelout<=1'b1;
23591: pixelout<=1'b1;
23592: pixelout<=1'b1;
23593: pixelout<=1'b1;
23594: pixelout<=1'b1;
23595: pixelout<=1'b1;
23596: pixelout<=1'b1;
23597: pixelout<=1'b1;
23598: pixelout<=1'b1;
23599: pixelout<=1'b1;
23600: pixelout<=1'b1;
23601: pixelout<=1'b1;
23602: pixelout<=1'b1;
23603: pixelout<=1'b1;
23604: pixelout<=1'b1;
23605: pixelout<=1'b1;
23606: pixelout<=1'b1;
23607: pixelout<=1'b1;
23608: pixelout<=1'b1;
23609: pixelout<=1'b1;
23610: pixelout<=1'b1;
23611: pixelout<=1'b1;
23612: pixelout<=1'b1;
23613: pixelout<=1'b1;
23614: pixelout<=1'b1;
23615: pixelout<=1'b1;
23616: pixelout<=1'b1;
23617: pixelout<=1'b1;
23618: pixelout<=1'b1;
23619: pixelout<=1'b1;
23620: pixelout<=1'b0;
23621: pixelout<=1'b0;
23622: pixelout<=1'b1;
23623: pixelout<=1'b0;
23624: pixelout<=1'b1;
23625: pixelout<=1'b0;
23626: pixelout<=1'b0;
23627: pixelout<=1'b0;
23628: pixelout<=1'b0;
23629: pixelout<=1'b1;
23630: pixelout<=1'b1;
23631: pixelout<=1'b1;
23632: pixelout<=1'b1;
23633: pixelout<=1'b1;
23634: pixelout<=1'b1;
23635: pixelout<=1'b1;
23636: pixelout<=1'b1;
23637: pixelout<=1'b1;
23638: pixelout<=1'b0;
23639: pixelout<=1'b1;
23640: pixelout<=1'b1;
23641: pixelout<=1'b1;
23642: pixelout<=1'b1;
23643: pixelout<=1'b0;
23644: pixelout<=1'b0;
23645: pixelout<=1'b0;
23646: pixelout<=1'b1;
23647: pixelout<=1'b1;
23648: pixelout<=1'b1;
23649: pixelout<=1'b0;
23650: pixelout<=1'b0;
23651: pixelout<=1'b0;
23652: pixelout<=1'b1;
23653: pixelout<=1'b1;
23654: pixelout<=1'b1;
23655: pixelout<=1'b1;
23656: pixelout<=1'b0;
23657: pixelout<=1'b0;
23658: pixelout<=1'b0;
23659: pixelout<=1'b1;
23660: pixelout<=1'b1;
23661: pixelout<=1'b0;
23662: pixelout<=1'b1;
23663: pixelout<=1'b1;
23664: pixelout<=1'b1;
23665: pixelout<=1'b1;
23666: pixelout<=1'b1;
23667: pixelout<=1'b1;
23668: pixelout<=1'b1;
23669: pixelout<=1'b1;
23670: pixelout<=1'b1;
23671: pixelout<=1'b1;
23672: pixelout<=1'b1;
23673: pixelout<=1'b1;
23674: pixelout<=1'b1;
23675: pixelout<=1'b1;
23676: pixelout<=1'b1;
23677: pixelout<=1'b1;
23678: pixelout<=1'b1;
23679: pixelout<=1'b1;
23680: pixelout<=1'b1;
23681: pixelout<=1'b1;
23682: pixelout<=1'b1;
23683: pixelout<=1'b1;
23684: pixelout<=1'b1;
23685: pixelout<=1'b1;
23686: pixelout<=1'b1;
23687: pixelout<=1'b1;
23688: pixelout<=1'b1;
23689: pixelout<=1'b1;
23690: pixelout<=1'b1;
23691: pixelout<=1'b1;
23692: pixelout<=1'b1;
23693: pixelout<=1'b1;
23694: pixelout<=1'b1;
23695: pixelout<=1'b1;
23696: pixelout<=1'b1;
23697: pixelout<=1'b1;
23698: pixelout<=1'b1;
23699: pixelout<=1'b1;
23700: pixelout<=1'b1;
23701: pixelout<=1'b1;
23702: pixelout<=1'b1;
23703: pixelout<=1'b1;
23704: pixelout<=1'b1;
23705: pixelout<=1'b1;
23706: pixelout<=1'b1;
23707: pixelout<=1'b1;
23708: pixelout<=1'b1;
23709: pixelout<=1'b1;
23710: pixelout<=1'b1;
23711: pixelout<=1'b1;
23712: pixelout<=1'b1;
23713: pixelout<=1'b1;
23714: pixelout<=1'b1;
23715: pixelout<=1'b1;
23716: pixelout<=1'b1;
23717: pixelout<=1'b1;
23718: pixelout<=1'b1;
23719: pixelout<=1'b1;
23720: pixelout<=1'b1;
23721: pixelout<=1'b1;
23722: pixelout<=1'b1;
23723: pixelout<=1'b1;
23724: pixelout<=1'b1;
23725: pixelout<=1'b1;
23726: pixelout<=1'b1;
23727: pixelout<=1'b1;
23728: pixelout<=1'b1;
23729: pixelout<=1'b1;
23730: pixelout<=1'b1;
23731: pixelout<=1'b1;
23732: pixelout<=1'b1;
23733: pixelout<=1'b1;
23734: pixelout<=1'b1;
23735: pixelout<=1'b1;
23736: pixelout<=1'b1;
23737: pixelout<=1'b1;
23738: pixelout<=1'b1;
23739: pixelout<=1'b1;
23740: pixelout<=1'b1;
23741: pixelout<=1'b1;
23742: pixelout<=1'b1;
23743: pixelout<=1'b1;
23744: pixelout<=1'b1;
23745: pixelout<=1'b1;
23746: pixelout<=1'b1;
23747: pixelout<=1'b1;
23748: pixelout<=1'b1;
23749: pixelout<=1'b1;
23750: pixelout<=1'b1;
23751: pixelout<=1'b1;
23752: pixelout<=1'b1;
23753: pixelout<=1'b1;
23754: pixelout<=1'b1;
23755: pixelout<=1'b1;
23756: pixelout<=1'b1;
23757: pixelout<=1'b1;
23758: pixelout<=1'b1;
23759: pixelout<=1'b1;
23760: pixelout<=1'b1;
23761: pixelout<=1'b1;
23762: pixelout<=1'b1;
23763: pixelout<=1'b1;
23764: pixelout<=1'b1;
23765: pixelout<=1'b1;
23766: pixelout<=1'b1;
23767: pixelout<=1'b1;
23768: pixelout<=1'b1;
23769: pixelout<=1'b1;
23770: pixelout<=1'b1;
23771: pixelout<=1'b1;
23772: pixelout<=1'b1;
23773: pixelout<=1'b1;
23774: pixelout<=1'b1;
23775: pixelout<=1'b1;
23776: pixelout<=1'b1;
23777: pixelout<=1'b1;
23778: pixelout<=1'b1;
23779: pixelout<=1'b1;
23780: pixelout<=1'b1;
23781: pixelout<=1'b1;
23782: pixelout<=1'b1;
23783: pixelout<=1'b1;
23784: pixelout<=1'b1;
23785: pixelout<=1'b1;
23786: pixelout<=1'b1;
23787: pixelout<=1'b1;
23788: pixelout<=1'b1;
23789: pixelout<=1'b1;
23790: pixelout<=1'b1;
23791: pixelout<=1'b1;
23792: pixelout<=1'b1;
23793: pixelout<=1'b1;
23794: pixelout<=1'b1;
23795: pixelout<=1'b1;
23796: pixelout<=1'b1;
23797: pixelout<=1'b1;
23798: pixelout<=1'b1;
23799: pixelout<=1'b1;
23800: pixelout<=1'b1;
23801: pixelout<=1'b1;
23802: pixelout<=1'b1;
23803: pixelout<=1'b1;
23804: pixelout<=1'b1;
23805: pixelout<=1'b1;
23806: pixelout<=1'b1;
23807: pixelout<=1'b1;
23808: pixelout<=1'b1;
23809: pixelout<=1'b1;
23810: pixelout<=1'b1;
23811: pixelout<=1'b1;
23812: pixelout<=1'b1;
23813: pixelout<=1'b1;
23814: pixelout<=1'b1;
23815: pixelout<=1'b1;
23816: pixelout<=1'b1;
23817: pixelout<=1'b1;
23818: pixelout<=1'b1;
23819: pixelout<=1'b1;
23820: pixelout<=1'b1;
23821: pixelout<=1'b1;
23822: pixelout<=1'b1;
23823: pixelout<=1'b1;
23824: pixelout<=1'b1;
23825: pixelout<=1'b1;
23826: pixelout<=1'b1;
23827: pixelout<=1'b1;
23828: pixelout<=1'b1;
23829: pixelout<=1'b1;
23830: pixelout<=1'b1;
23831: pixelout<=1'b1;
23832: pixelout<=1'b1;
23833: pixelout<=1'b1;
23834: pixelout<=1'b1;
23835: pixelout<=1'b1;
23836: pixelout<=1'b1;
23837: pixelout<=1'b1;
23838: pixelout<=1'b1;
23839: pixelout<=1'b1;
23840: pixelout<=1'b1;
23841: pixelout<=1'b1;
23842: pixelout<=1'b1;
23843: pixelout<=1'b1;
23844: pixelout<=1'b1;
23845: pixelout<=1'b1;
23846: pixelout<=1'b1;
23847: pixelout<=1'b1;
23848: pixelout<=1'b1;
23849: pixelout<=1'b1;
23850: pixelout<=1'b1;
23851: pixelout<=1'b1;
23852: pixelout<=1'b1;
23853: pixelout<=1'b1;
23854: pixelout<=1'b1;
23855: pixelout<=1'b1;
23856: pixelout<=1'b1;
23857: pixelout<=1'b1;
23858: pixelout<=1'b1;
23859: pixelout<=1'b1;
23860: pixelout<=1'b1;
23861: pixelout<=1'b1;
23862: pixelout<=1'b1;
23863: pixelout<=1'b1;
23864: pixelout<=1'b1;
23865: pixelout<=1'b1;
23866: pixelout<=1'b1;
23867: pixelout<=1'b1;
23868: pixelout<=1'b1;
23869: pixelout<=1'b1;
23870: pixelout<=1'b1;
23871: pixelout<=1'b1;
23872: pixelout<=1'b1;
23873: pixelout<=1'b1;
23874: pixelout<=1'b1;
23875: pixelout<=1'b1;
23876: pixelout<=1'b1;
23877: pixelout<=1'b1;
23878: pixelout<=1'b1;
23879: pixelout<=1'b1;
23880: pixelout<=1'b1;
23881: pixelout<=1'b1;
23882: pixelout<=1'b1;
23883: pixelout<=1'b1;
23884: pixelout<=1'b1;
23885: pixelout<=1'b1;
23886: pixelout<=1'b1;
23887: pixelout<=1'b1;
23888: pixelout<=1'b1;
23889: pixelout<=1'b1;
23890: pixelout<=1'b1;
23891: pixelout<=1'b1;
23892: pixelout<=1'b1;
23893: pixelout<=1'b1;
23894: pixelout<=1'b1;
23895: pixelout<=1'b1;
23896: pixelout<=1'b1;
23897: pixelout<=1'b1;
23898: pixelout<=1'b1;
23899: pixelout<=1'b1;
23900: pixelout<=1'b1;
23901: pixelout<=1'b1;
23902: pixelout<=1'b1;
23903: pixelout<=1'b1;
23904: pixelout<=1'b1;
23905: pixelout<=1'b1;
23906: pixelout<=1'b1;
23907: pixelout<=1'b1;
23908: pixelout<=1'b1;
23909: pixelout<=1'b1;
23910: pixelout<=1'b1;
23911: pixelout<=1'b1;
23912: pixelout<=1'b1;
23913: pixelout<=1'b1;
23914: pixelout<=1'b1;
23915: pixelout<=1'b1;
23916: pixelout<=1'b1;
23917: pixelout<=1'b1;
23918: pixelout<=1'b1;
23919: pixelout<=1'b1;
23920: pixelout<=1'b1;
23921: pixelout<=1'b1;
23922: pixelout<=1'b1;
23923: pixelout<=1'b1;
23924: pixelout<=1'b1;
23925: pixelout<=1'b1;
23926: pixelout<=1'b1;
23927: pixelout<=1'b1;
23928: pixelout<=1'b1;
23929: pixelout<=1'b1;
23930: pixelout<=1'b1;
23931: pixelout<=1'b1;
23932: pixelout<=1'b1;
23933: pixelout<=1'b1;
23934: pixelout<=1'b1;
23935: pixelout<=1'b1;
23936: pixelout<=1'b1;
23937: pixelout<=1'b1;
23938: pixelout<=1'b1;
23939: pixelout<=1'b1;
23940: pixelout<=1'b1;
23941: pixelout<=1'b1;
23942: pixelout<=1'b1;
23943: pixelout<=1'b1;
23944: pixelout<=1'b1;
23945: pixelout<=1'b1;
23946: pixelout<=1'b1;
23947: pixelout<=1'b1;
23948: pixelout<=1'b1;
23949: pixelout<=1'b1;
23950: pixelout<=1'b1;
23951: pixelout<=1'b1;
23952: pixelout<=1'b1;
23953: pixelout<=1'b1;
23954: pixelout<=1'b1;
23955: pixelout<=1'b1;
23956: pixelout<=1'b1;
23957: pixelout<=1'b1;
23958: pixelout<=1'b1;
23959: pixelout<=1'b1;
23960: pixelout<=1'b1;
23961: pixelout<=1'b1;
23962: pixelout<=1'b1;
23963: pixelout<=1'b1;
23964: pixelout<=1'b1;
23965: pixelout<=1'b1;
23966: pixelout<=1'b1;
23967: pixelout<=1'b1;
23968: pixelout<=1'b1;
23969: pixelout<=1'b1;
23970: pixelout<=1'b1;
23971: pixelout<=1'b1;
23972: pixelout<=1'b1;
23973: pixelout<=1'b1;
23974: pixelout<=1'b1;
23975: pixelout<=1'b1;
23976: pixelout<=1'b1;
23977: pixelout<=1'b1;
23978: pixelout<=1'b1;
23979: pixelout<=1'b1;
23980: pixelout<=1'b1;
23981: pixelout<=1'b1;
23982: pixelout<=1'b1;
23983: pixelout<=1'b1;
23984: pixelout<=1'b1;
23985: pixelout<=1'b1;
23986: pixelout<=1'b1;
23987: pixelout<=1'b1;
23988: pixelout<=1'b1;
23989: pixelout<=1'b1;
23990: pixelout<=1'b1;
23991: pixelout<=1'b1;
23992: pixelout<=1'b1;
23993: pixelout<=1'b1;
23994: pixelout<=1'b1;
23995: pixelout<=1'b1;
23996: pixelout<=1'b1;
23997: pixelout<=1'b1;
23998: pixelout<=1'b1;
23999: pixelout<=1'b1;
24000: pixelout<=1'b1;
24001: pixelout<=1'b1;
24002: pixelout<=1'b1;
24003: pixelout<=1'b1;
24004: pixelout<=1'b1;
24005: pixelout<=1'b1;
24006: pixelout<=1'b1;
24007: pixelout<=1'b1;
24008: pixelout<=1'b1;
24009: pixelout<=1'b1;
24010: pixelout<=1'b1;
24011: pixelout<=1'b1;
24012: pixelout<=1'b1;
24013: pixelout<=1'b1;
24014: pixelout<=1'b1;
24015: pixelout<=1'b1;
24016: pixelout<=1'b1;
24017: pixelout<=1'b1;
24018: pixelout<=1'b1;
24019: pixelout<=1'b1;
24020: pixelout<=1'b1;
24021: pixelout<=1'b1;
24022: pixelout<=1'b1;
24023: pixelout<=1'b1;
24024: pixelout<=1'b1;
24025: pixelout<=1'b1;
24026: pixelout<=1'b1;
24027: pixelout<=1'b1;
24028: pixelout<=1'b1;
24029: pixelout<=1'b1;
24030: pixelout<=1'b1;
24031: pixelout<=1'b1;
24032: pixelout<=1'b1;
24033: pixelout<=1'b1;
24034: pixelout<=1'b1;
24035: pixelout<=1'b1;
24036: pixelout<=1'b1;
24037: pixelout<=1'b1;
24038: pixelout<=1'b1;
24039: pixelout<=1'b1;
24040: pixelout<=1'b1;
24041: pixelout<=1'b1;
24042: pixelout<=1'b1;
24043: pixelout<=1'b1;
24044: pixelout<=1'b1;
24045: pixelout<=1'b1;
24046: pixelout<=1'b1;
24047: pixelout<=1'b1;
24048: pixelout<=1'b1;
24049: pixelout<=1'b1;
24050: pixelout<=1'b1;
24051: pixelout<=1'b1;
24052: pixelout<=1'b1;
24053: pixelout<=1'b1;
24054: pixelout<=1'b1;
24055: pixelout<=1'b1;
24056: pixelout<=1'b1;
24057: pixelout<=1'b1;
24058: pixelout<=1'b1;
24059: pixelout<=1'b1;
24060: pixelout<=1'b1;
24061: pixelout<=1'b1;
24062: pixelout<=1'b1;
24063: pixelout<=1'b1;
24064: pixelout<=1'b1;
24065: pixelout<=1'b1;
24066: pixelout<=1'b1;
24067: pixelout<=1'b1;
24068: pixelout<=1'b1;
24069: pixelout<=1'b1;
24070: pixelout<=1'b1;
24071: pixelout<=1'b1;
24072: pixelout<=1'b1;
24073: pixelout<=1'b1;
24074: pixelout<=1'b1;
24075: pixelout<=1'b1;
24076: pixelout<=1'b1;
24077: pixelout<=1'b1;
24078: pixelout<=1'b1;
24079: pixelout<=1'b1;
24080: pixelout<=1'b1;
24081: pixelout<=1'b1;
24082: pixelout<=1'b1;
24083: pixelout<=1'b1;
24084: pixelout<=1'b1;
24085: pixelout<=1'b1;
24086: pixelout<=1'b1;
24087: pixelout<=1'b1;
24088: pixelout<=1'b1;
24089: pixelout<=1'b1;
24090: pixelout<=1'b1;
24091: pixelout<=1'b1;
24092: pixelout<=1'b1;
24093: pixelout<=1'b1;
24094: pixelout<=1'b1;
24095: pixelout<=1'b1;
24096: pixelout<=1'b1;
24097: pixelout<=1'b1;
24098: pixelout<=1'b1;
24099: pixelout<=1'b1;
24100: pixelout<=1'b1;
24101: pixelout<=1'b1;
24102: pixelout<=1'b1;
24103: pixelout<=1'b1;
24104: pixelout<=1'b1;
24105: pixelout<=1'b1;
24106: pixelout<=1'b1;
24107: pixelout<=1'b1;
24108: pixelout<=1'b1;
24109: pixelout<=1'b1;
24110: pixelout<=1'b1;
24111: pixelout<=1'b1;
24112: pixelout<=1'b1;
24113: pixelout<=1'b1;
24114: pixelout<=1'b1;
24115: pixelout<=1'b1;
24116: pixelout<=1'b1;
24117: pixelout<=1'b1;
24118: pixelout<=1'b1;
24119: pixelout<=1'b1;
24120: pixelout<=1'b1;
24121: pixelout<=1'b1;
24122: pixelout<=1'b1;
24123: pixelout<=1'b1;
24124: pixelout<=1'b1;
24125: pixelout<=1'b1;
24126: pixelout<=1'b1;
24127: pixelout<=1'b1;
24128: pixelout<=1'b1;
24129: pixelout<=1'b1;
24130: pixelout<=1'b1;
24131: pixelout<=1'b1;
24132: pixelout<=1'b1;
24133: pixelout<=1'b1;
24134: pixelout<=1'b1;
24135: pixelout<=1'b1;
24136: pixelout<=1'b1;
24137: pixelout<=1'b1;
24138: pixelout<=1'b1;
24139: pixelout<=1'b1;
24140: pixelout<=1'b1;
24141: pixelout<=1'b1;
24142: pixelout<=1'b1;
24143: pixelout<=1'b1;
24144: pixelout<=1'b1;
24145: pixelout<=1'b1;
24146: pixelout<=1'b1;
24147: pixelout<=1'b1;
24148: pixelout<=1'b1;
24149: pixelout<=1'b1;
24150: pixelout<=1'b1;
24151: pixelout<=1'b1;
24152: pixelout<=1'b1;
24153: pixelout<=1'b1;
24154: pixelout<=1'b1;
24155: pixelout<=1'b1;
24156: pixelout<=1'b1;
24157: pixelout<=1'b1;
24158: pixelout<=1'b1;
24159: pixelout<=1'b1;
24160: pixelout<=1'b1;
24161: pixelout<=1'b1;
24162: pixelout<=1'b1;
24163: pixelout<=1'b1;
24164: pixelout<=1'b1;
24165: pixelout<=1'b1;
24166: pixelout<=1'b1;
24167: pixelout<=1'b1;
24168: pixelout<=1'b1;
24169: pixelout<=1'b1;
24170: pixelout<=1'b1;
24171: pixelout<=1'b1;
24172: pixelout<=1'b1;
24173: pixelout<=1'b1;
24174: pixelout<=1'b1;
24175: pixelout<=1'b1;
24176: pixelout<=1'b1;
24177: pixelout<=1'b1;
24178: pixelout<=1'b1;
24179: pixelout<=1'b1;
24180: pixelout<=1'b1;
24181: pixelout<=1'b1;
24182: pixelout<=1'b1;
24183: pixelout<=1'b1;
24184: pixelout<=1'b1;
24185: pixelout<=1'b1;
24186: pixelout<=1'b1;
24187: pixelout<=1'b1;
24188: pixelout<=1'b1;
24189: pixelout<=1'b1;
24190: pixelout<=1'b1;
24191: pixelout<=1'b1;
24192: pixelout<=1'b1;
24193: pixelout<=1'b1;
24194: pixelout<=1'b1;
24195: pixelout<=1'b1;
24196: pixelout<=1'b1;
24197: pixelout<=1'b1;
24198: pixelout<=1'b1;
24199: pixelout<=1'b1;
24200: pixelout<=1'b1;
24201: pixelout<=1'b1;
24202: pixelout<=1'b1;
24203: pixelout<=1'b1;
24204: pixelout<=1'b1;
24205: pixelout<=1'b1;
24206: pixelout<=1'b1;
24207: pixelout<=1'b1;
24208: pixelout<=1'b1;
24209: pixelout<=1'b1;
24210: pixelout<=1'b1;
24211: pixelout<=1'b1;
24212: pixelout<=1'b1;
24213: pixelout<=1'b1;
24214: pixelout<=1'b1;
24215: pixelout<=1'b1;
24216: pixelout<=1'b1;
24217: pixelout<=1'b1;
24218: pixelout<=1'b1;
24219: pixelout<=1'b1;
24220: pixelout<=1'b1;
24221: pixelout<=1'b1;
24222: pixelout<=1'b1;
24223: pixelout<=1'b1;
24224: pixelout<=1'b1;
24225: pixelout<=1'b1;
24226: pixelout<=1'b1;
24227: pixelout<=1'b1;
24228: pixelout<=1'b1;
24229: pixelout<=1'b1;
24230: pixelout<=1'b1;
24231: pixelout<=1'b1;
24232: pixelout<=1'b1;
24233: pixelout<=1'b1;
24234: pixelout<=1'b1;
24235: pixelout<=1'b1;
24236: pixelout<=1'b1;
24237: pixelout<=1'b1;
24238: pixelout<=1'b1;
24239: pixelout<=1'b1;
24240: pixelout<=1'b1;
24241: pixelout<=1'b1;
24242: pixelout<=1'b1;
24243: pixelout<=1'b1;
24244: pixelout<=1'b1;
24245: pixelout<=1'b1;
24246: pixelout<=1'b1;
24247: pixelout<=1'b1;
24248: pixelout<=1'b1;
24249: pixelout<=1'b1;
24250: pixelout<=1'b1;
24251: pixelout<=1'b1;
24252: pixelout<=1'b1;
24253: pixelout<=1'b1;
24254: pixelout<=1'b1;
24255: pixelout<=1'b1;
24256: pixelout<=1'b1;
24257: pixelout<=1'b1;
24258: pixelout<=1'b1;
24259: pixelout<=1'b1;
24260: pixelout<=1'b1;
24261: pixelout<=1'b1;
24262: pixelout<=1'b1;
24263: pixelout<=1'b1;
24264: pixelout<=1'b1;
24265: pixelout<=1'b1;
24266: pixelout<=1'b1;
24267: pixelout<=1'b1;
24268: pixelout<=1'b1;
24269: pixelout<=1'b1;
24270: pixelout<=1'b1;
24271: pixelout<=1'b1;
24272: pixelout<=1'b1;
24273: pixelout<=1'b1;
24274: pixelout<=1'b1;
24275: pixelout<=1'b1;
24276: pixelout<=1'b1;
24277: pixelout<=1'b1;
24278: pixelout<=1'b1;
24279: pixelout<=1'b1;
24280: pixelout<=1'b1;
24281: pixelout<=1'b1;
24282: pixelout<=1'b1;
24283: pixelout<=1'b1;
24284: pixelout<=1'b1;
24285: pixelout<=1'b1;
24286: pixelout<=1'b1;
24287: pixelout<=1'b1;
24288: pixelout<=1'b1;
24289: pixelout<=1'b1;
24290: pixelout<=1'b1;
24291: pixelout<=1'b1;
24292: pixelout<=1'b1;
24293: pixelout<=1'b1;
24294: pixelout<=1'b1;
24295: pixelout<=1'b1;
24296: pixelout<=1'b1;
24297: pixelout<=1'b1;
24298: pixelout<=1'b1;
24299: pixelout<=1'b1;
24300: pixelout<=1'b1;
24301: pixelout<=1'b1;
24302: pixelout<=1'b1;
24303: pixelout<=1'b1;
24304: pixelout<=1'b1;
24305: pixelout<=1'b1;
24306: pixelout<=1'b1;
24307: pixelout<=1'b1;
24308: pixelout<=1'b1;
24309: pixelout<=1'b1;
24310: pixelout<=1'b1;
24311: pixelout<=1'b1;
24312: pixelout<=1'b1;
24313: pixelout<=1'b1;
24314: pixelout<=1'b1;
24315: pixelout<=1'b1;
24316: pixelout<=1'b1;
24317: pixelout<=1'b1;
24318: pixelout<=1'b1;
24319: pixelout<=1'b1;
24320: pixelout<=1'b1;
24321: pixelout<=1'b1;
24322: pixelout<=1'b1;
24323: pixelout<=1'b1;
24324: pixelout<=1'b1;
24325: pixelout<=1'b1;
24326: pixelout<=1'b1;
24327: pixelout<=1'b1;
24328: pixelout<=1'b1;
24329: pixelout<=1'b1;
24330: pixelout<=1'b1;
24331: pixelout<=1'b1;
24332: pixelout<=1'b1;
24333: pixelout<=1'b1;
24334: pixelout<=1'b1;
24335: pixelout<=1'b1;
24336: pixelout<=1'b1;
24337: pixelout<=1'b1;
24338: pixelout<=1'b1;
24339: pixelout<=1'b1;
24340: pixelout<=1'b1;
24341: pixelout<=1'b1;
24342: pixelout<=1'b1;
24343: pixelout<=1'b1;
24344: pixelout<=1'b1;
24345: pixelout<=1'b1;
24346: pixelout<=1'b1;
24347: pixelout<=1'b1;
24348: pixelout<=1'b1;
24349: pixelout<=1'b1;
24350: pixelout<=1'b1;
24351: pixelout<=1'b1;
24352: pixelout<=1'b1;
24353: pixelout<=1'b1;
24354: pixelout<=1'b1;
24355: pixelout<=1'b1;
24356: pixelout<=1'b1;
24357: pixelout<=1'b1;
24358: pixelout<=1'b1;
24359: pixelout<=1'b1;
24360: pixelout<=1'b1;
24361: pixelout<=1'b1;
24362: pixelout<=1'b1;
24363: pixelout<=1'b1;
24364: pixelout<=1'b1;
24365: pixelout<=1'b1;
24366: pixelout<=1'b1;
24367: pixelout<=1'b1;
24368: pixelout<=1'b1;
24369: pixelout<=1'b1;
24370: pixelout<=1'b1;
24371: pixelout<=1'b1;
24372: pixelout<=1'b1;
24373: pixelout<=1'b1;
24374: pixelout<=1'b1;
24375: pixelout<=1'b1;
24376: pixelout<=1'b1;
24377: pixelout<=1'b1;
24378: pixelout<=1'b1;
24379: pixelout<=1'b1;
24380: pixelout<=1'b1;
24381: pixelout<=1'b1;
24382: pixelout<=1'b1;
24383: pixelout<=1'b1;
24384: pixelout<=1'b1;
24385: pixelout<=1'b1;
24386: pixelout<=1'b1;
24387: pixelout<=1'b1;
24388: pixelout<=1'b1;
24389: pixelout<=1'b1;
24390: pixelout<=1'b1;
24391: pixelout<=1'b1;
24392: pixelout<=1'b1;
24393: pixelout<=1'b1;
24394: pixelout<=1'b1;
24395: pixelout<=1'b1;
24396: pixelout<=1'b1;
24397: pixelout<=1'b1;
24398: pixelout<=1'b1;
24399: pixelout<=1'b1;
24400: pixelout<=1'b1;
24401: pixelout<=1'b1;
24402: pixelout<=1'b1;
24403: pixelout<=1'b1;
24404: pixelout<=1'b1;
24405: pixelout<=1'b1;
24406: pixelout<=1'b1;
24407: pixelout<=1'b1;
24408: pixelout<=1'b1;
24409: pixelout<=1'b1;
24410: pixelout<=1'b1;
24411: pixelout<=1'b1;
24412: pixelout<=1'b1;
24413: pixelout<=1'b1;
24414: pixelout<=1'b1;
24415: pixelout<=1'b1;
24416: pixelout<=1'b1;
24417: pixelout<=1'b1;
24418: pixelout<=1'b1;
24419: pixelout<=1'b1;
24420: pixelout<=1'b1;
24421: pixelout<=1'b1;
24422: pixelout<=1'b1;
24423: pixelout<=1'b1;
24424: pixelout<=1'b1;
24425: pixelout<=1'b1;
24426: pixelout<=1'b1;
24427: pixelout<=1'b1;
24428: pixelout<=1'b1;
24429: pixelout<=1'b1;
24430: pixelout<=1'b1;
24431: pixelout<=1'b1;
24432: pixelout<=1'b1;
24433: pixelout<=1'b1;
24434: pixelout<=1'b1;
24435: pixelout<=1'b1;
24436: pixelout<=1'b1;
24437: pixelout<=1'b1;
24438: pixelout<=1'b1;
24439: pixelout<=1'b1;
24440: pixelout<=1'b1;
24441: pixelout<=1'b1;
24442: pixelout<=1'b1;
24443: pixelout<=1'b1;
24444: pixelout<=1'b1;
24445: pixelout<=1'b1;
24446: pixelout<=1'b1;
24447: pixelout<=1'b1;
24448: pixelout<=1'b1;
24449: pixelout<=1'b1;
24450: pixelout<=1'b1;
24451: pixelout<=1'b1;
24452: pixelout<=1'b1;
24453: pixelout<=1'b1;
24454: pixelout<=1'b1;
24455: pixelout<=1'b1;
24456: pixelout<=1'b1;
24457: pixelout<=1'b1;
24458: pixelout<=1'b1;
24459: pixelout<=1'b1;
24460: pixelout<=1'b1;
24461: pixelout<=1'b1;
24462: pixelout<=1'b1;
24463: pixelout<=1'b1;
24464: pixelout<=1'b1;
24465: pixelout<=1'b1;
24466: pixelout<=1'b1;
24467: pixelout<=1'b1;
24468: pixelout<=1'b1;
24469: pixelout<=1'b1;
24470: pixelout<=1'b1;
24471: pixelout<=1'b1;
24472: pixelout<=1'b1;
24473: pixelout<=1'b1;
24474: pixelout<=1'b1;
24475: pixelout<=1'b1;
24476: pixelout<=1'b1;
24477: pixelout<=1'b1;
24478: pixelout<=1'b1;
24479: pixelout<=1'b1;
24480: pixelout<=1'b1;
24481: pixelout<=1'b1;
24482: pixelout<=1'b1;
24483: pixelout<=1'b1;
24484: pixelout<=1'b1;
24485: pixelout<=1'b1;
24486: pixelout<=1'b1;
24487: pixelout<=1'b1;
24488: pixelout<=1'b1;
24489: pixelout<=1'b1;
24490: pixelout<=1'b1;
24491: pixelout<=1'b1;
24492: pixelout<=1'b1;
24493: pixelout<=1'b1;
24494: pixelout<=1'b1;
24495: pixelout<=1'b1;
24496: pixelout<=1'b1;
24497: pixelout<=1'b1;
24498: pixelout<=1'b1;
24499: pixelout<=1'b1;
24500: pixelout<=1'b1;
24501: pixelout<=1'b1;
24502: pixelout<=1'b1;
24503: pixelout<=1'b1;
24504: pixelout<=1'b1;
24505: pixelout<=1'b1;
24506: pixelout<=1'b1;
24507: pixelout<=1'b1;
24508: pixelout<=1'b1;
24509: pixelout<=1'b1;
24510: pixelout<=1'b1;
24511: pixelout<=1'b1;
24512: pixelout<=1'b1;
24513: pixelout<=1'b1;
24514: pixelout<=1'b1;
24515: pixelout<=1'b1;
24516: pixelout<=1'b1;
24517: pixelout<=1'b1;
24518: pixelout<=1'b1;
24519: pixelout<=1'b1;
24520: pixelout<=1'b1;
24521: pixelout<=1'b1;
24522: pixelout<=1'b1;
24523: pixelout<=1'b1;
24524: pixelout<=1'b1;
24525: pixelout<=1'b1;
24526: pixelout<=1'b1;
24527: pixelout<=1'b1;
24528: pixelout<=1'b1;
24529: pixelout<=1'b1;
24530: pixelout<=1'b1;
24531: pixelout<=1'b1;
24532: pixelout<=1'b1;
24533: pixelout<=1'b1;
24534: pixelout<=1'b1;
24535: pixelout<=1'b1;
24536: pixelout<=1'b1;
24537: pixelout<=1'b1;
24538: pixelout<=1'b1;
24539: pixelout<=1'b1;
24540: pixelout<=1'b1;
24541: pixelout<=1'b1;
24542: pixelout<=1'b1;
24543: pixelout<=1'b1;
24544: pixelout<=1'b1;
24545: pixelout<=1'b1;
24546: pixelout<=1'b1;
24547: pixelout<=1'b1;
24548: pixelout<=1'b1;
24549: pixelout<=1'b1;
24550: pixelout<=1'b1;
24551: pixelout<=1'b1;
24552: pixelout<=1'b1;
24553: pixelout<=1'b1;
24554: pixelout<=1'b1;
24555: pixelout<=1'b1;
24556: pixelout<=1'b1;
24557: pixelout<=1'b1;
24558: pixelout<=1'b1;
24559: pixelout<=1'b1;
24560: pixelout<=1'b1;
24561: pixelout<=1'b1;
24562: pixelout<=1'b1;
24563: pixelout<=1'b1;
24564: pixelout<=1'b1;
24565: pixelout<=1'b1;
24566: pixelout<=1'b1;
24567: pixelout<=1'b1;
24568: pixelout<=1'b1;
24569: pixelout<=1'b1;
24570: pixelout<=1'b1;
24571: pixelout<=1'b1;
24572: pixelout<=1'b1;
24573: pixelout<=1'b1;
24574: pixelout<=1'b1;
24575: pixelout<=1'b1;
24576: pixelout<=1'b1;
24577: pixelout<=1'b1;
24578: pixelout<=1'b1;
24579: pixelout<=1'b1;
24580: pixelout<=1'b1;
24581: pixelout<=1'b1;
24582: pixelout<=1'b1;
24583: pixelout<=1'b1;
24584: pixelout<=1'b1;
24585: pixelout<=1'b1;
24586: pixelout<=1'b1;
24587: pixelout<=1'b1;
24588: pixelout<=1'b1;
24589: pixelout<=1'b1;
24590: pixelout<=1'b1;
24591: pixelout<=1'b1;
24592: pixelout<=1'b1;
24593: pixelout<=1'b1;
24594: pixelout<=1'b1;
24595: pixelout<=1'b1;
24596: pixelout<=1'b1;
24597: pixelout<=1'b1;
24598: pixelout<=1'b1;
24599: pixelout<=1'b1;
24600: pixelout<=1'b1;
24601: pixelout<=1'b1;
24602: pixelout<=1'b1;
24603: pixelout<=1'b1;
24604: pixelout<=1'b1;
24605: pixelout<=1'b1;
24606: pixelout<=1'b1;
24607: pixelout<=1'b1;
24608: pixelout<=1'b1;
24609: pixelout<=1'b1;
24610: pixelout<=1'b1;
24611: pixelout<=1'b1;
24612: pixelout<=1'b1;
24613: pixelout<=1'b1;
24614: pixelout<=1'b1;
24615: pixelout<=1'b1;
24616: pixelout<=1'b1;
24617: pixelout<=1'b1;
24618: pixelout<=1'b1;
24619: pixelout<=1'b1;
24620: pixelout<=1'b1;
24621: pixelout<=1'b1;
24622: pixelout<=1'b1;
24623: pixelout<=1'b1;
24624: pixelout<=1'b1;
24625: pixelout<=1'b1;
24626: pixelout<=1'b1;
24627: pixelout<=1'b1;
24628: pixelout<=1'b1;
24629: pixelout<=1'b1;
24630: pixelout<=1'b1;
24631: pixelout<=1'b1;
24632: pixelout<=1'b1;
24633: pixelout<=1'b1;
24634: pixelout<=1'b1;
24635: pixelout<=1'b1;
24636: pixelout<=1'b1;
24637: pixelout<=1'b1;
24638: pixelout<=1'b1;
24639: pixelout<=1'b1;
24640: pixelout<=1'b1;
24641: pixelout<=1'b1;
24642: pixelout<=1'b1;
24643: pixelout<=1'b1;
24644: pixelout<=1'b1;
24645: pixelout<=1'b1;
24646: pixelout<=1'b1;
24647: pixelout<=1'b1;
24648: pixelout<=1'b1;
24649: pixelout<=1'b1;
24650: pixelout<=1'b1;
24651: pixelout<=1'b1;
24652: pixelout<=1'b1;
24653: pixelout<=1'b1;
24654: pixelout<=1'b1;
24655: pixelout<=1'b1;
24656: pixelout<=1'b1;
24657: pixelout<=1'b1;
24658: pixelout<=1'b1;
24659: pixelout<=1'b1;
24660: pixelout<=1'b1;
24661: pixelout<=1'b1;
24662: pixelout<=1'b1;
24663: pixelout<=1'b1;
24664: pixelout<=1'b1;
24665: pixelout<=1'b1;
24666: pixelout<=1'b1;
24667: pixelout<=1'b1;
24668: pixelout<=1'b1;
24669: pixelout<=1'b1;
24670: pixelout<=1'b1;
24671: pixelout<=1'b1;
24672: pixelout<=1'b1;
24673: pixelout<=1'b1;
24674: pixelout<=1'b1;
24675: pixelout<=1'b1;
24676: pixelout<=1'b1;
24677: pixelout<=1'b1;
24678: pixelout<=1'b1;
24679: pixelout<=1'b1;
24680: pixelout<=1'b1;
24681: pixelout<=1'b1;
24682: pixelout<=1'b1;
24683: pixelout<=1'b1;
24684: pixelout<=1'b1;
24685: pixelout<=1'b1;
24686: pixelout<=1'b1;
24687: pixelout<=1'b1;
24688: pixelout<=1'b1;
24689: pixelout<=1'b1;
24690: pixelout<=1'b1;
24691: pixelout<=1'b1;
24692: pixelout<=1'b1;
24693: pixelout<=1'b1;
24694: pixelout<=1'b1;
24695: pixelout<=1'b1;
24696: pixelout<=1'b1;
24697: pixelout<=1'b1;
24698: pixelout<=1'b1;
24699: pixelout<=1'b1;
24700: pixelout<=1'b1;
24701: pixelout<=1'b1;
24702: pixelout<=1'b1;
24703: pixelout<=1'b1;
24704: pixelout<=1'b1;
24705: pixelout<=1'b1;
24706: pixelout<=1'b1;
24707: pixelout<=1'b1;
24708: pixelout<=1'b1;
24709: pixelout<=1'b1;
24710: pixelout<=1'b1;
24711: pixelout<=1'b1;
24712: pixelout<=1'b1;
24713: pixelout<=1'b1;
24714: pixelout<=1'b1;
24715: pixelout<=1'b1;
24716: pixelout<=1'b1;
24717: pixelout<=1'b1;
24718: pixelout<=1'b1;
24719: pixelout<=1'b1;
24720: pixelout<=1'b1;
24721: pixelout<=1'b1;
24722: pixelout<=1'b1;
24723: pixelout<=1'b1;
24724: pixelout<=1'b1;
24725: pixelout<=1'b1;
24726: pixelout<=1'b1;
24727: pixelout<=1'b1;
24728: pixelout<=1'b1;
24729: pixelout<=1'b1;
24730: pixelout<=1'b1;
24731: pixelout<=1'b1;
24732: pixelout<=1'b1;
24733: pixelout<=1'b1;
24734: pixelout<=1'b1;
24735: pixelout<=1'b1;
24736: pixelout<=1'b1;
24737: pixelout<=1'b1;
24738: pixelout<=1'b1;
24739: pixelout<=1'b1;
24740: pixelout<=1'b1;
24741: pixelout<=1'b1;
24742: pixelout<=1'b1;
24743: pixelout<=1'b1;
24744: pixelout<=1'b1;
24745: pixelout<=1'b1;
24746: pixelout<=1'b1;
24747: pixelout<=1'b1;
24748: pixelout<=1'b1;
24749: pixelout<=1'b1;
24750: pixelout<=1'b1;
24751: pixelout<=1'b1;
24752: pixelout<=1'b1;
24753: pixelout<=1'b1;
24754: pixelout<=1'b1;
24755: pixelout<=1'b1;
24756: pixelout<=1'b1;
24757: pixelout<=1'b1;
24758: pixelout<=1'b1;
24759: pixelout<=1'b1;
24760: pixelout<=1'b1;
24761: pixelout<=1'b1;
24762: pixelout<=1'b1;
24763: pixelout<=1'b1;
24764: pixelout<=1'b1;
24765: pixelout<=1'b1;
24766: pixelout<=1'b1;
24767: pixelout<=1'b1;
24768: pixelout<=1'b1;
24769: pixelout<=1'b1;
24770: pixelout<=1'b1;
24771: pixelout<=1'b1;
24772: pixelout<=1'b1;
24773: pixelout<=1'b1;
24774: pixelout<=1'b1;
24775: pixelout<=1'b1;
24776: pixelout<=1'b1;
24777: pixelout<=1'b1;
24778: pixelout<=1'b1;
24779: pixelout<=1'b1;
24780: pixelout<=1'b1;
24781: pixelout<=1'b1;
24782: pixelout<=1'b1;
24783: pixelout<=1'b1;
24784: pixelout<=1'b1;
24785: pixelout<=1'b1;
24786: pixelout<=1'b1;
24787: pixelout<=1'b1;
24788: pixelout<=1'b1;
24789: pixelout<=1'b1;
24790: pixelout<=1'b1;
24791: pixelout<=1'b1;
24792: pixelout<=1'b1;
24793: pixelout<=1'b1;
24794: pixelout<=1'b1;
24795: pixelout<=1'b1;
24796: pixelout<=1'b1;
24797: pixelout<=1'b1;
24798: pixelout<=1'b1;
24799: pixelout<=1'b1;
24800: pixelout<=1'b1;
24801: pixelout<=1'b1;
24802: pixelout<=1'b1;
24803: pixelout<=1'b1;
24804: pixelout<=1'b1;
24805: pixelout<=1'b1;
24806: pixelout<=1'b1;
24807: pixelout<=1'b1;
24808: pixelout<=1'b1;
24809: pixelout<=1'b1;
24810: pixelout<=1'b1;
24811: pixelout<=1'b1;
24812: pixelout<=1'b1;
24813: pixelout<=1'b1;
24814: pixelout<=1'b1;
24815: pixelout<=1'b1;
24816: pixelout<=1'b1;
24817: pixelout<=1'b1;
24818: pixelout<=1'b1;
24819: pixelout<=1'b1;
24820: pixelout<=1'b1;
24821: pixelout<=1'b1;
24822: pixelout<=1'b1;
24823: pixelout<=1'b1;
24824: pixelout<=1'b1;
24825: pixelout<=1'b1;
24826: pixelout<=1'b1;
24827: pixelout<=1'b1;
24828: pixelout<=1'b1;
24829: pixelout<=1'b1;
24830: pixelout<=1'b1;
24831: pixelout<=1'b1;
24832: pixelout<=1'b1;
24833: pixelout<=1'b1;
24834: pixelout<=1'b1;
24835: pixelout<=1'b1;
24836: pixelout<=1'b1;
24837: pixelout<=1'b1;
24838: pixelout<=1'b1;
24839: pixelout<=1'b1;
24840: pixelout<=1'b1;
24841: pixelout<=1'b1;
24842: pixelout<=1'b1;
24843: pixelout<=1'b1;
24844: pixelout<=1'b1;
24845: pixelout<=1'b1;
24846: pixelout<=1'b1;
24847: pixelout<=1'b1;
24848: pixelout<=1'b1;
24849: pixelout<=1'b1;
24850: pixelout<=1'b1;
24851: pixelout<=1'b1;
24852: pixelout<=1'b1;
24853: pixelout<=1'b1;
24854: pixelout<=1'b1;
24855: pixelout<=1'b1;
24856: pixelout<=1'b1;
24857: pixelout<=1'b1;
24858: pixelout<=1'b1;
24859: pixelout<=1'b1;
24860: pixelout<=1'b1;
24861: pixelout<=1'b1;
24862: pixelout<=1'b1;
24863: pixelout<=1'b1;
24864: pixelout<=1'b1;
24865: pixelout<=1'b1;
24866: pixelout<=1'b1;
24867: pixelout<=1'b1;
24868: pixelout<=1'b1;
24869: pixelout<=1'b1;
24870: pixelout<=1'b1;
24871: pixelout<=1'b1;
24872: pixelout<=1'b1;
24873: pixelout<=1'b1;
24874: pixelout<=1'b1;
24875: pixelout<=1'b1;
24876: pixelout<=1'b1;
24877: pixelout<=1'b1;
24878: pixelout<=1'b1;
24879: pixelout<=1'b1;
24880: pixelout<=1'b1;
24881: pixelout<=1'b1;
24882: pixelout<=1'b1;
24883: pixelout<=1'b1;
24884: pixelout<=1'b1;
24885: pixelout<=1'b1;
24886: pixelout<=1'b1;
24887: pixelout<=1'b1;
24888: pixelout<=1'b1;
24889: pixelout<=1'b1;
24890: pixelout<=1'b1;
24891: pixelout<=1'b1;
24892: pixelout<=1'b1;
24893: pixelout<=1'b1;
24894: pixelout<=1'b1;
24895: pixelout<=1'b1;
24896: pixelout<=1'b1;
24897: pixelout<=1'b1;
24898: pixelout<=1'b1;
24899: pixelout<=1'b1;
24900: pixelout<=1'b1;
24901: pixelout<=1'b1;
24902: pixelout<=1'b1;
24903: pixelout<=1'b1;
24904: pixelout<=1'b1;
24905: pixelout<=1'b1;
24906: pixelout<=1'b1;
24907: pixelout<=1'b1;
24908: pixelout<=1'b1;
24909: pixelout<=1'b1;
24910: pixelout<=1'b1;
24911: pixelout<=1'b1;
24912: pixelout<=1'b1;
24913: pixelout<=1'b1;
24914: pixelout<=1'b1;
24915: pixelout<=1'b1;
24916: pixelout<=1'b1;
24917: pixelout<=1'b1;
24918: pixelout<=1'b1;
24919: pixelout<=1'b1;
24920: pixelout<=1'b1;
24921: pixelout<=1'b1;
24922: pixelout<=1'b1;
24923: pixelout<=1'b1;
24924: pixelout<=1'b1;
24925: pixelout<=1'b1;
24926: pixelout<=1'b1;
24927: pixelout<=1'b1;
24928: pixelout<=1'b1;
24929: pixelout<=1'b1;
24930: pixelout<=1'b1;
24931: pixelout<=1'b1;
24932: pixelout<=1'b1;
24933: pixelout<=1'b1;
24934: pixelout<=1'b1;
24935: pixelout<=1'b1;
24936: pixelout<=1'b1;
24937: pixelout<=1'b1;
24938: pixelout<=1'b1;
24939: pixelout<=1'b1;
24940: pixelout<=1'b1;
24941: pixelout<=1'b1;
24942: pixelout<=1'b1;
24943: pixelout<=1'b1;
24944: pixelout<=1'b1;
24945: pixelout<=1'b1;
24946: pixelout<=1'b1;
24947: pixelout<=1'b1;
24948: pixelout<=1'b1;
24949: pixelout<=1'b1;
24950: pixelout<=1'b1;
24951: pixelout<=1'b1;
24952: pixelout<=1'b1;
24953: pixelout<=1'b1;
24954: pixelout<=1'b1;
24955: pixelout<=1'b1;
24956: pixelout<=1'b1;
24957: pixelout<=1'b1;
24958: pixelout<=1'b1;
24959: pixelout<=1'b1;
24960: pixelout<=1'b1;
24961: pixelout<=1'b1;
24962: pixelout<=1'b1;
24963: pixelout<=1'b1;
24964: pixelout<=1'b1;
24965: pixelout<=1'b1;
24966: pixelout<=1'b1;
24967: pixelout<=1'b1;
24968: pixelout<=1'b1;
24969: pixelout<=1'b1;
24970: pixelout<=1'b1;
24971: pixelout<=1'b1;
24972: pixelout<=1'b1;
24973: pixelout<=1'b1;
24974: pixelout<=1'b1;
24975: pixelout<=1'b1;
24976: pixelout<=1'b1;
24977: pixelout<=1'b1;
24978: pixelout<=1'b1;
24979: pixelout<=1'b1;
24980: pixelout<=1'b1;
24981: pixelout<=1'b1;
24982: pixelout<=1'b1;
24983: pixelout<=1'b1;
24984: pixelout<=1'b1;
24985: pixelout<=1'b1;
24986: pixelout<=1'b1;
24987: pixelout<=1'b1;
24988: pixelout<=1'b1;
24989: pixelout<=1'b1;
24990: pixelout<=1'b1;
24991: pixelout<=1'b1;
24992: pixelout<=1'b1;
24993: pixelout<=1'b1;
24994: pixelout<=1'b1;
24995: pixelout<=1'b1;
24996: pixelout<=1'b1;
24997: pixelout<=1'b1;
24998: pixelout<=1'b1;
24999: pixelout<=1'b1;
25000: pixelout<=1'b1;
25001: pixelout<=1'b1;
25002: pixelout<=1'b1;
25003: pixelout<=1'b1;
25004: pixelout<=1'b1;
25005: pixelout<=1'b1;
25006: pixelout<=1'b1;
25007: pixelout<=1'b1;
25008: pixelout<=1'b1;
25009: pixelout<=1'b1;
25010: pixelout<=1'b1;
25011: pixelout<=1'b1;
25012: pixelout<=1'b1;
25013: pixelout<=1'b1;
25014: pixelout<=1'b1;
25015: pixelout<=1'b1;
25016: pixelout<=1'b1;
25017: pixelout<=1'b1;
25018: pixelout<=1'b1;
25019: pixelout<=1'b1;
25020: pixelout<=1'b1;
25021: pixelout<=1'b1;
25022: pixelout<=1'b1;
25023: pixelout<=1'b1;
25024: pixelout<=1'b1;
25025: pixelout<=1'b1;
25026: pixelout<=1'b1;
25027: pixelout<=1'b1;
25028: pixelout<=1'b1;
25029: pixelout<=1'b1;
25030: pixelout<=1'b1;
25031: pixelout<=1'b1;
25032: pixelout<=1'b1;
25033: pixelout<=1'b1;
25034: pixelout<=1'b1;
25035: pixelout<=1'b1;
25036: pixelout<=1'b1;
25037: pixelout<=1'b1;
25038: pixelout<=1'b1;
25039: pixelout<=1'b1;
25040: pixelout<=1'b1;
25041: pixelout<=1'b1;
25042: pixelout<=1'b1;
25043: pixelout<=1'b1;
25044: pixelout<=1'b1;
25045: pixelout<=1'b1;
25046: pixelout<=1'b1;
25047: pixelout<=1'b1;
25048: pixelout<=1'b1;
25049: pixelout<=1'b1;
25050: pixelout<=1'b1;
25051: pixelout<=1'b1;
25052: pixelout<=1'b1;
25053: pixelout<=1'b1;
25054: pixelout<=1'b1;
25055: pixelout<=1'b1;
25056: pixelout<=1'b1;
25057: pixelout<=1'b1;
25058: pixelout<=1'b1;
25059: pixelout<=1'b1;
25060: pixelout<=1'b1;
25061: pixelout<=1'b1;
25062: pixelout<=1'b1;
25063: pixelout<=1'b1;
25064: pixelout<=1'b1;
25065: pixelout<=1'b1;
25066: pixelout<=1'b1;
25067: pixelout<=1'b1;
25068: pixelout<=1'b1;
25069: pixelout<=1'b1;
25070: pixelout<=1'b1;
25071: pixelout<=1'b1;
25072: pixelout<=1'b1;
25073: pixelout<=1'b1;
25074: pixelout<=1'b1;
25075: pixelout<=1'b1;
25076: pixelout<=1'b1;
25077: pixelout<=1'b1;
25078: pixelout<=1'b1;
25079: pixelout<=1'b1;
25080: pixelout<=1'b1;
25081: pixelout<=1'b1;
25082: pixelout<=1'b1;
25083: pixelout<=1'b1;
25084: pixelout<=1'b1;
25085: pixelout<=1'b1;
25086: pixelout<=1'b1;
25087: pixelout<=1'b1;
25088: pixelout<=1'b1;
25089: pixelout<=1'b1;
25090: pixelout<=1'b1;
25091: pixelout<=1'b1;
25092: pixelout<=1'b1;
25093: pixelout<=1'b1;
25094: pixelout<=1'b1;
25095: pixelout<=1'b1;
25096: pixelout<=1'b1;
25097: pixelout<=1'b1;
25098: pixelout<=1'b1;
25099: pixelout<=1'b1;
25100: pixelout<=1'b1;
25101: pixelout<=1'b1;
25102: pixelout<=1'b1;
25103: pixelout<=1'b1;
25104: pixelout<=1'b1;
25105: pixelout<=1'b1;
25106: pixelout<=1'b1;
25107: pixelout<=1'b1;
25108: pixelout<=1'b1;
25109: pixelout<=1'b1;
25110: pixelout<=1'b1;
25111: pixelout<=1'b1;
25112: pixelout<=1'b1;
25113: pixelout<=1'b1;
25114: pixelout<=1'b1;
25115: pixelout<=1'b1;
25116: pixelout<=1'b1;
25117: pixelout<=1'b1;
25118: pixelout<=1'b1;
25119: pixelout<=1'b1;
25120: pixelout<=1'b1;
25121: pixelout<=1'b1;
25122: pixelout<=1'b1;
25123: pixelout<=1'b1;
25124: pixelout<=1'b1;
25125: pixelout<=1'b1;
25126: pixelout<=1'b1;
25127: pixelout<=1'b1;
25128: pixelout<=1'b1;
25129: pixelout<=1'b1;
25130: pixelout<=1'b1;
25131: pixelout<=1'b1;
25132: pixelout<=1'b1;
25133: pixelout<=1'b1;
25134: pixelout<=1'b1;
25135: pixelout<=1'b1;
25136: pixelout<=1'b1;
25137: pixelout<=1'b1;
25138: pixelout<=1'b1;
25139: pixelout<=1'b1;
25140: pixelout<=1'b1;
25141: pixelout<=1'b1;
25142: pixelout<=1'b1;
25143: pixelout<=1'b1;
25144: pixelout<=1'b1;
25145: pixelout<=1'b1;
25146: pixelout<=1'b1;
25147: pixelout<=1'b1;
25148: pixelout<=1'b1;
25149: pixelout<=1'b1;
25150: pixelout<=1'b1;
25151: pixelout<=1'b1;
25152: pixelout<=1'b1;
25153: pixelout<=1'b1;
25154: pixelout<=1'b1;
25155: pixelout<=1'b1;
25156: pixelout<=1'b1;
25157: pixelout<=1'b1;
25158: pixelout<=1'b1;
25159: pixelout<=1'b1;
25160: pixelout<=1'b1;
25161: pixelout<=1'b1;
25162: pixelout<=1'b1;
25163: pixelout<=1'b1;
25164: pixelout<=1'b1;
25165: pixelout<=1'b1;
25166: pixelout<=1'b1;
25167: pixelout<=1'b1;
25168: pixelout<=1'b1;
25169: pixelout<=1'b1;
25170: pixelout<=1'b1;
25171: pixelout<=1'b1;
25172: pixelout<=1'b1;
25173: pixelout<=1'b1;
25174: pixelout<=1'b1;
25175: pixelout<=1'b1;
25176: pixelout<=1'b1;
25177: pixelout<=1'b1;
25178: pixelout<=1'b1;
25179: pixelout<=1'b1;
25180: pixelout<=1'b1;
25181: pixelout<=1'b1;
25182: pixelout<=1'b1;
25183: pixelout<=1'b1;
25184: pixelout<=1'b1;
25185: pixelout<=1'b1;
25186: pixelout<=1'b1;
25187: pixelout<=1'b1;
25188: pixelout<=1'b1;
25189: pixelout<=1'b1;
25190: pixelout<=1'b1;
25191: pixelout<=1'b1;
25192: pixelout<=1'b1;
25193: pixelout<=1'b1;
25194: pixelout<=1'b1;
25195: pixelout<=1'b1;
25196: pixelout<=1'b1;
25197: pixelout<=1'b1;
25198: pixelout<=1'b1;
25199: pixelout<=1'b1;
25200: pixelout<=1'b1;
25201: pixelout<=1'b1;
25202: pixelout<=1'b1;
25203: pixelout<=1'b1;
25204: pixelout<=1'b1;
25205: pixelout<=1'b1;
25206: pixelout<=1'b1;
25207: pixelout<=1'b1;
25208: pixelout<=1'b1;
25209: pixelout<=1'b1;
25210: pixelout<=1'b1;
25211: pixelout<=1'b1;
25212: pixelout<=1'b1;
25213: pixelout<=1'b1;
25214: pixelout<=1'b1;
25215: pixelout<=1'b1;
25216: pixelout<=1'b1;
25217: pixelout<=1'b1;
25218: pixelout<=1'b1;
25219: pixelout<=1'b1;
25220: pixelout<=1'b1;
25221: pixelout<=1'b1;
25222: pixelout<=1'b1;
25223: pixelout<=1'b1;
25224: pixelout<=1'b1;
25225: pixelout<=1'b1;
25226: pixelout<=1'b1;
25227: pixelout<=1'b1;
25228: pixelout<=1'b1;
25229: pixelout<=1'b1;
25230: pixelout<=1'b1;
25231: pixelout<=1'b1;
25232: pixelout<=1'b1;
25233: pixelout<=1'b1;
25234: pixelout<=1'b1;
25235: pixelout<=1'b1;
25236: pixelout<=1'b1;
25237: pixelout<=1'b1;
25238: pixelout<=1'b1;
25239: pixelout<=1'b1;
25240: pixelout<=1'b1;
25241: pixelout<=1'b1;
25242: pixelout<=1'b1;
25243: pixelout<=1'b1;
25244: pixelout<=1'b1;
25245: pixelout<=1'b1;
25246: pixelout<=1'b1;
25247: pixelout<=1'b1;
25248: pixelout<=1'b1;
25249: pixelout<=1'b1;
25250: pixelout<=1'b1;
25251: pixelout<=1'b1;
25252: pixelout<=1'b1;
25253: pixelout<=1'b1;
25254: pixelout<=1'b1;
25255: pixelout<=1'b1;
25256: pixelout<=1'b1;
25257: pixelout<=1'b1;
25258: pixelout<=1'b1;
25259: pixelout<=1'b1;
25260: pixelout<=1'b1;
25261: pixelout<=1'b1;
25262: pixelout<=1'b1;
25263: pixelout<=1'b1;
25264: pixelout<=1'b1;
25265: pixelout<=1'b1;
25266: pixelout<=1'b1;
25267: pixelout<=1'b1;
25268: pixelout<=1'b1;
25269: pixelout<=1'b1;
25270: pixelout<=1'b1;
25271: pixelout<=1'b1;
25272: pixelout<=1'b1;
25273: pixelout<=1'b1;
25274: pixelout<=1'b1;
25275: pixelout<=1'b1;
25276: pixelout<=1'b1;
25277: pixelout<=1'b1;
25278: pixelout<=1'b1;
25279: pixelout<=1'b1;
25280: pixelout<=1'b1;
25281: pixelout<=1'b1;
25282: pixelout<=1'b1;
25283: pixelout<=1'b1;
25284: pixelout<=1'b1;
25285: pixelout<=1'b1;
25286: pixelout<=1'b1;
25287: pixelout<=1'b1;
25288: pixelout<=1'b1;
25289: pixelout<=1'b1;
25290: pixelout<=1'b1;
25291: pixelout<=1'b1;
25292: pixelout<=1'b1;
25293: pixelout<=1'b1;
25294: pixelout<=1'b1;
25295: pixelout<=1'b1;
25296: pixelout<=1'b1;
25297: pixelout<=1'b1;
25298: pixelout<=1'b1;
25299: pixelout<=1'b1;
25300: pixelout<=1'b1;
25301: pixelout<=1'b1;
25302: pixelout<=1'b1;
25303: pixelout<=1'b1;
25304: pixelout<=1'b1;
25305: pixelout<=1'b1;
25306: pixelout<=1'b1;
25307: pixelout<=1'b1;
25308: pixelout<=1'b1;
25309: pixelout<=1'b1;
25310: pixelout<=1'b1;
25311: pixelout<=1'b1;
25312: pixelout<=1'b1;
25313: pixelout<=1'b1;
25314: pixelout<=1'b1;
25315: pixelout<=1'b1;
25316: pixelout<=1'b1;
25317: pixelout<=1'b1;
25318: pixelout<=1'b1;
25319: pixelout<=1'b1;
25320: pixelout<=1'b1;
25321: pixelout<=1'b1;
25322: pixelout<=1'b1;
25323: pixelout<=1'b1;
25324: pixelout<=1'b1;
25325: pixelout<=1'b1;
25326: pixelout<=1'b1;
25327: pixelout<=1'b1;
25328: pixelout<=1'b1;
25329: pixelout<=1'b1;
25330: pixelout<=1'b1;
25331: pixelout<=1'b1;
25332: pixelout<=1'b1;
25333: pixelout<=1'b1;
25334: pixelout<=1'b1;
25335: pixelout<=1'b1;
25336: pixelout<=1'b1;
25337: pixelout<=1'b1;
25338: pixelout<=1'b1;
25339: pixelout<=1'b1;
25340: pixelout<=1'b1;
25341: pixelout<=1'b1;
25342: pixelout<=1'b1;
25343: pixelout<=1'b1;
25344: pixelout<=1'b1;
25345: pixelout<=1'b1;
25346: pixelout<=1'b1;
25347: pixelout<=1'b1;
25348: pixelout<=1'b1;
25349: pixelout<=1'b1;
25350: pixelout<=1'b1;
25351: pixelout<=1'b1;
25352: pixelout<=1'b1;
25353: pixelout<=1'b1;
25354: pixelout<=1'b1;
25355: pixelout<=1'b1;
25356: pixelout<=1'b1;
25357: pixelout<=1'b1;
25358: pixelout<=1'b1;
25359: pixelout<=1'b1;
25360: pixelout<=1'b1;
25361: pixelout<=1'b1;
25362: pixelout<=1'b1;
25363: pixelout<=1'b1;
25364: pixelout<=1'b1;
25365: pixelout<=1'b1;
25366: pixelout<=1'b1;
25367: pixelout<=1'b1;
25368: pixelout<=1'b1;
25369: pixelout<=1'b1;
25370: pixelout<=1'b1;
25371: pixelout<=1'b1;
25372: pixelout<=1'b1;
25373: pixelout<=1'b1;
25374: pixelout<=1'b1;
25375: pixelout<=1'b1;
25376: pixelout<=1'b1;
25377: pixelout<=1'b1;
25378: pixelout<=1'b1;
25379: pixelout<=1'b1;
25380: pixelout<=1'b1;
25381: pixelout<=1'b1;
25382: pixelout<=1'b1;
25383: pixelout<=1'b1;
25384: pixelout<=1'b1;
25385: pixelout<=1'b1;
25386: pixelout<=1'b1;
25387: pixelout<=1'b1;
25388: pixelout<=1'b1;
25389: pixelout<=1'b1;
25390: pixelout<=1'b1;
25391: pixelout<=1'b1;
25392: pixelout<=1'b1;
25393: pixelout<=1'b1;
25394: pixelout<=1'b1;
25395: pixelout<=1'b1;
25396: pixelout<=1'b1;
25397: pixelout<=1'b1;
25398: pixelout<=1'b1;
25399: pixelout<=1'b1;
25400: pixelout<=1'b1;
25401: pixelout<=1'b1;
25402: pixelout<=1'b1;
25403: pixelout<=1'b1;
25404: pixelout<=1'b1;
25405: pixelout<=1'b1;
25406: pixelout<=1'b1;
25407: pixelout<=1'b1;
25408: pixelout<=1'b1;
25409: pixelout<=1'b1;
25410: pixelout<=1'b1;
25411: pixelout<=1'b1;
25412: pixelout<=1'b1;
25413: pixelout<=1'b1;
25414: pixelout<=1'b1;
25415: pixelout<=1'b1;
25416: pixelout<=1'b1;
25417: pixelout<=1'b1;
25418: pixelout<=1'b1;
25419: pixelout<=1'b1;
25420: pixelout<=1'b1;
25421: pixelout<=1'b1;
25422: pixelout<=1'b1;
25423: pixelout<=1'b1;
25424: pixelout<=1'b1;
25425: pixelout<=1'b1;
25426: pixelout<=1'b1;
25427: pixelout<=1'b1;
25428: pixelout<=1'b1;
25429: pixelout<=1'b1;
25430: pixelout<=1'b1;
25431: pixelout<=1'b1;
25432: pixelout<=1'b1;
25433: pixelout<=1'b1;
25434: pixelout<=1'b1;
25435: pixelout<=1'b1;
25436: pixelout<=1'b1;
25437: pixelout<=1'b1;
25438: pixelout<=1'b1;
25439: pixelout<=1'b1;
25440: pixelout<=1'b1;
25441: pixelout<=1'b1;
25442: pixelout<=1'b1;
25443: pixelout<=1'b1;
25444: pixelout<=1'b1;
25445: pixelout<=1'b1;
25446: pixelout<=1'b1;
25447: pixelout<=1'b1;
25448: pixelout<=1'b1;
25449: pixelout<=1'b1;
25450: pixelout<=1'b1;
25451: pixelout<=1'b1;
25452: pixelout<=1'b1;
25453: pixelout<=1'b1;
25454: pixelout<=1'b1;
25455: pixelout<=1'b1;
25456: pixelout<=1'b1;
25457: pixelout<=1'b1;
25458: pixelout<=1'b1;
25459: pixelout<=1'b1;
25460: pixelout<=1'b1;
25461: pixelout<=1'b1;
25462: pixelout<=1'b1;
25463: pixelout<=1'b1;
25464: pixelout<=1'b1;
25465: pixelout<=1'b1;
25466: pixelout<=1'b1;
25467: pixelout<=1'b1;
25468: pixelout<=1'b1;
25469: pixelout<=1'b1;
25470: pixelout<=1'b1;
25471: pixelout<=1'b1;
25472: pixelout<=1'b1;
25473: pixelout<=1'b1;
25474: pixelout<=1'b1;
25475: pixelout<=1'b1;
25476: pixelout<=1'b1;
25477: pixelout<=1'b1;
25478: pixelout<=1'b1;
25479: pixelout<=1'b1;
25480: pixelout<=1'b1;
25481: pixelout<=1'b1;
25482: pixelout<=1'b1;
25483: pixelout<=1'b1;
25484: pixelout<=1'b1;
25485: pixelout<=1'b1;
25486: pixelout<=1'b1;
25487: pixelout<=1'b1;
25488: pixelout<=1'b1;
25489: pixelout<=1'b1;
25490: pixelout<=1'b1;
25491: pixelout<=1'b1;
25492: pixelout<=1'b1;
25493: pixelout<=1'b1;
25494: pixelout<=1'b1;
25495: pixelout<=1'b1;
25496: pixelout<=1'b1;
25497: pixelout<=1'b1;
25498: pixelout<=1'b1;
25499: pixelout<=1'b1;
25500: pixelout<=1'b1;
25501: pixelout<=1'b1;
25502: pixelout<=1'b1;
25503: pixelout<=1'b1;
25504: pixelout<=1'b1;
25505: pixelout<=1'b1;
25506: pixelout<=1'b1;
25507: pixelout<=1'b1;
25508: pixelout<=1'b1;
25509: pixelout<=1'b1;
25510: pixelout<=1'b1;
25511: pixelout<=1'b1;
25512: pixelout<=1'b1;
25513: pixelout<=1'b1;
25514: pixelout<=1'b1;
25515: pixelout<=1'b1;
25516: pixelout<=1'b1;
25517: pixelout<=1'b1;
25518: pixelout<=1'b1;
25519: pixelout<=1'b1;
25520: pixelout<=1'b1;
25521: pixelout<=1'b1;
25522: pixelout<=1'b1;
25523: pixelout<=1'b1;
25524: pixelout<=1'b1;
25525: pixelout<=1'b1;
25526: pixelout<=1'b1;
25527: pixelout<=1'b1;
25528: pixelout<=1'b1;
25529: pixelout<=1'b1;
25530: pixelout<=1'b1;
25531: pixelout<=1'b1;
25532: pixelout<=1'b1;
25533: pixelout<=1'b1;
25534: pixelout<=1'b1;
25535: pixelout<=1'b0;
25536: pixelout<=1'b0;
25537: pixelout<=1'b1;
25538: pixelout<=1'b1;
25539: pixelout<=1'b1;
25540: pixelout<=1'b1;
25541: pixelout<=1'b1;
25542: pixelout<=1'b1;
25543: pixelout<=1'b1;
25544: pixelout<=1'b1;
25545: pixelout<=1'b1;
25546: pixelout<=1'b1;
25547: pixelout<=1'b1;
25548: pixelout<=1'b1;
25549: pixelout<=1'b1;
25550: pixelout<=1'b1;
25551: pixelout<=1'b1;
25552: pixelout<=1'b1;
25553: pixelout<=1'b1;
25554: pixelout<=1'b1;
25555: pixelout<=1'b1;
25556: pixelout<=1'b1;
25557: pixelout<=1'b1;
25558: pixelout<=1'b1;
25559: pixelout<=1'b1;
25560: pixelout<=1'b1;
25561: pixelout<=1'b1;
25562: pixelout<=1'b1;
25563: pixelout<=1'b1;
25564: pixelout<=1'b1;
25565: pixelout<=1'b1;
25566: pixelout<=1'b1;
25567: pixelout<=1'b1;
25568: pixelout<=1'b1;
25569: pixelout<=1'b1;
25570: pixelout<=1'b1;
25571: pixelout<=1'b1;
25572: pixelout<=1'b1;
25573: pixelout<=1'b1;
25574: pixelout<=1'b1;
25575: pixelout<=1'b1;
25576: pixelout<=1'b1;
25577: pixelout<=1'b1;
25578: pixelout<=1'b1;
25579: pixelout<=1'b1;
25580: pixelout<=1'b1;
25581: pixelout<=1'b1;
25582: pixelout<=1'b1;
25583: pixelout<=1'b1;
25584: pixelout<=1'b1;
25585: pixelout<=1'b1;
25586: pixelout<=1'b1;
25587: pixelout<=1'b1;
25588: pixelout<=1'b1;
25589: pixelout<=1'b1;
25590: pixelout<=1'b1;
25591: pixelout<=1'b1;
25592: pixelout<=1'b1;
25593: pixelout<=1'b1;
25594: pixelout<=1'b1;
25595: pixelout<=1'b1;
25596: pixelout<=1'b1;
25597: pixelout<=1'b1;
25598: pixelout<=1'b1;
25599: pixelout<=1'b1;
25600: pixelout<=1'b1;
25601: pixelout<=1'b1;
25602: pixelout<=1'b1;
25603: pixelout<=1'b1;
25604: pixelout<=1'b1;
25605: pixelout<=1'b1;
25606: pixelout<=1'b1;
25607: pixelout<=1'b1;
25608: pixelout<=1'b1;
25609: pixelout<=1'b1;
25610: pixelout<=1'b1;
25611: pixelout<=1'b1;
25612: pixelout<=1'b1;
25613: pixelout<=1'b1;
25614: pixelout<=1'b1;
25615: pixelout<=1'b1;
25616: pixelout<=1'b1;
25617: pixelout<=1'b1;
25618: pixelout<=1'b1;
25619: pixelout<=1'b1;
25620: pixelout<=1'b1;
25621: pixelout<=1'b1;
25622: pixelout<=1'b1;
25623: pixelout<=1'b1;
25624: pixelout<=1'b1;
25625: pixelout<=1'b1;
25626: pixelout<=1'b1;
25627: pixelout<=1'b1;
25628: pixelout<=1'b1;
25629: pixelout<=1'b1;
25630: pixelout<=1'b1;
25631: pixelout<=1'b1;
25632: pixelout<=1'b1;
25633: pixelout<=1'b1;
25634: pixelout<=1'b1;
25635: pixelout<=1'b1;
25636: pixelout<=1'b1;
25637: pixelout<=1'b1;
25638: pixelout<=1'b1;
25639: pixelout<=1'b1;
25640: pixelout<=1'b1;
25641: pixelout<=1'b1;
25642: pixelout<=1'b1;
25643: pixelout<=1'b1;
25644: pixelout<=1'b1;
25645: pixelout<=1'b1;
25646: pixelout<=1'b1;
25647: pixelout<=1'b1;
25648: pixelout<=1'b1;
25649: pixelout<=1'b1;
25650: pixelout<=1'b1;
25651: pixelout<=1'b1;
25652: pixelout<=1'b1;
25653: pixelout<=1'b1;
25654: pixelout<=1'b1;
25655: pixelout<=1'b1;
25656: pixelout<=1'b1;
25657: pixelout<=1'b1;
25658: pixelout<=1'b1;
25659: pixelout<=1'b1;
25660: pixelout<=1'b1;
25661: pixelout<=1'b1;
25662: pixelout<=1'b1;
25663: pixelout<=1'b1;
25664: pixelout<=1'b1;
25665: pixelout<=1'b1;
25666: pixelout<=1'b1;
25667: pixelout<=1'b1;
25668: pixelout<=1'b1;
25669: pixelout<=1'b1;
25670: pixelout<=1'b1;
25671: pixelout<=1'b1;
25672: pixelout<=1'b1;
25673: pixelout<=1'b1;
25674: pixelout<=1'b1;
25675: pixelout<=1'b1;
25676: pixelout<=1'b1;
25677: pixelout<=1'b1;
25678: pixelout<=1'b1;
25679: pixelout<=1'b1;
25680: pixelout<=1'b1;
25681: pixelout<=1'b1;
25682: pixelout<=1'b1;
25683: pixelout<=1'b1;
25684: pixelout<=1'b1;
25685: pixelout<=1'b1;
25686: pixelout<=1'b1;
25687: pixelout<=1'b1;
25688: pixelout<=1'b1;
25689: pixelout<=1'b1;
25690: pixelout<=1'b1;
25691: pixelout<=1'b1;
25692: pixelout<=1'b1;
25693: pixelout<=1'b1;
25694: pixelout<=1'b1;
25695: pixelout<=1'b1;
25696: pixelout<=1'b1;
25697: pixelout<=1'b1;
25698: pixelout<=1'b1;
25699: pixelout<=1'b1;
25700: pixelout<=1'b1;
25701: pixelout<=1'b1;
25702: pixelout<=1'b1;
25703: pixelout<=1'b1;
25704: pixelout<=1'b1;
25705: pixelout<=1'b1;
25706: pixelout<=1'b1;
25707: pixelout<=1'b1;
25708: pixelout<=1'b1;
25709: pixelout<=1'b1;
25710: pixelout<=1'b1;
25711: pixelout<=1'b1;
25712: pixelout<=1'b1;
25713: pixelout<=1'b1;
25714: pixelout<=1'b1;
25715: pixelout<=1'b1;
25716: pixelout<=1'b1;
25717: pixelout<=1'b1;
25718: pixelout<=1'b1;
25719: pixelout<=1'b1;
25720: pixelout<=1'b1;
25721: pixelout<=1'b1;
25722: pixelout<=1'b1;
25723: pixelout<=1'b1;
25724: pixelout<=1'b1;
25725: pixelout<=1'b1;
25726: pixelout<=1'b1;
25727: pixelout<=1'b1;
25728: pixelout<=1'b1;
25729: pixelout<=1'b1;
25730: pixelout<=1'b1;
25731: pixelout<=1'b1;
25732: pixelout<=1'b1;
25733: pixelout<=1'b1;
25734: pixelout<=1'b1;
25735: pixelout<=1'b1;
25736: pixelout<=1'b1;
25737: pixelout<=1'b1;
25738: pixelout<=1'b1;
25739: pixelout<=1'b1;
25740: pixelout<=1'b1;
25741: pixelout<=1'b1;
25742: pixelout<=1'b1;
25743: pixelout<=1'b1;
25744: pixelout<=1'b1;
25745: pixelout<=1'b1;
25746: pixelout<=1'b1;
25747: pixelout<=1'b1;
25748: pixelout<=1'b1;
25749: pixelout<=1'b1;
25750: pixelout<=1'b1;
25751: pixelout<=1'b1;
25752: pixelout<=1'b1;
25753: pixelout<=1'b1;
25754: pixelout<=1'b1;
25755: pixelout<=1'b1;
25756: pixelout<=1'b1;
25757: pixelout<=1'b1;
25758: pixelout<=1'b1;
25759: pixelout<=1'b1;
25760: pixelout<=1'b1;
25761: pixelout<=1'b1;
25762: pixelout<=1'b1;
25763: pixelout<=1'b1;
25764: pixelout<=1'b1;
25765: pixelout<=1'b1;
25766: pixelout<=1'b1;
25767: pixelout<=1'b1;
25768: pixelout<=1'b1;
25769: pixelout<=1'b1;
25770: pixelout<=1'b1;
25771: pixelout<=1'b1;
25772: pixelout<=1'b1;
25773: pixelout<=1'b1;
25774: pixelout<=1'b1;
25775: pixelout<=1'b1;
25776: pixelout<=1'b0;
25777: pixelout<=1'b1;
25778: pixelout<=1'b1;
25779: pixelout<=1'b1;
25780: pixelout<=1'b1;
25781: pixelout<=1'b1;
25782: pixelout<=1'b1;
25783: pixelout<=1'b1;
25784: pixelout<=1'b1;
25785: pixelout<=1'b1;
25786: pixelout<=1'b1;
25787: pixelout<=1'b1;
25788: pixelout<=1'b1;
25789: pixelout<=1'b1;
25790: pixelout<=1'b1;
25791: pixelout<=1'b1;
25792: pixelout<=1'b1;
25793: pixelout<=1'b1;
25794: pixelout<=1'b1;
25795: pixelout<=1'b1;
25796: pixelout<=1'b1;
25797: pixelout<=1'b1;
25798: pixelout<=1'b1;
25799: pixelout<=1'b1;
25800: pixelout<=1'b1;
25801: pixelout<=1'b1;
25802: pixelout<=1'b1;
25803: pixelout<=1'b1;
25804: pixelout<=1'b1;
25805: pixelout<=1'b1;
25806: pixelout<=1'b1;
25807: pixelout<=1'b1;
25808: pixelout<=1'b1;
25809: pixelout<=1'b1;
25810: pixelout<=1'b1;
25811: pixelout<=1'b1;
25812: pixelout<=1'b1;
25813: pixelout<=1'b1;
25814: pixelout<=1'b1;
25815: pixelout<=1'b1;
25816: pixelout<=1'b1;
25817: pixelout<=1'b1;
25818: pixelout<=1'b1;
25819: pixelout<=1'b1;
25820: pixelout<=1'b1;
25821: pixelout<=1'b1;
25822: pixelout<=1'b1;
25823: pixelout<=1'b1;
25824: pixelout<=1'b1;
25825: pixelout<=1'b1;
25826: pixelout<=1'b1;
25827: pixelout<=1'b1;
25828: pixelout<=1'b1;
25829: pixelout<=1'b1;
25830: pixelout<=1'b1;
25831: pixelout<=1'b1;
25832: pixelout<=1'b1;
25833: pixelout<=1'b1;
25834: pixelout<=1'b1;
25835: pixelout<=1'b1;
25836: pixelout<=1'b1;
25837: pixelout<=1'b1;
25838: pixelout<=1'b1;
25839: pixelout<=1'b1;
25840: pixelout<=1'b1;
25841: pixelout<=1'b1;
25842: pixelout<=1'b1;
25843: pixelout<=1'b1;
25844: pixelout<=1'b1;
25845: pixelout<=1'b1;
25846: pixelout<=1'b1;
25847: pixelout<=1'b1;
25848: pixelout<=1'b1;
25849: pixelout<=1'b1;
25850: pixelout<=1'b1;
25851: pixelout<=1'b1;
25852: pixelout<=1'b1;
25853: pixelout<=1'b1;
25854: pixelout<=1'b1;
25855: pixelout<=1'b1;
25856: pixelout<=1'b1;
25857: pixelout<=1'b1;
25858: pixelout<=1'b1;
25859: pixelout<=1'b1;
25860: pixelout<=1'b1;
25861: pixelout<=1'b1;
25862: pixelout<=1'b1;
25863: pixelout<=1'b1;
25864: pixelout<=1'b1;
25865: pixelout<=1'b1;
25866: pixelout<=1'b1;
25867: pixelout<=1'b1;
25868: pixelout<=1'b1;
25869: pixelout<=1'b1;
25870: pixelout<=1'b1;
25871: pixelout<=1'b1;
25872: pixelout<=1'b1;
25873: pixelout<=1'b1;
25874: pixelout<=1'b1;
25875: pixelout<=1'b1;
25876: pixelout<=1'b1;
25877: pixelout<=1'b1;
25878: pixelout<=1'b1;
25879: pixelout<=1'b1;
25880: pixelout<=1'b1;
25881: pixelout<=1'b1;
25882: pixelout<=1'b1;
25883: pixelout<=1'b1;
25884: pixelout<=1'b1;
25885: pixelout<=1'b1;
25886: pixelout<=1'b1;
25887: pixelout<=1'b1;
25888: pixelout<=1'b1;
25889: pixelout<=1'b1;
25890: pixelout<=1'b1;
25891: pixelout<=1'b1;
25892: pixelout<=1'b1;
25893: pixelout<=1'b1;
25894: pixelout<=1'b1;
25895: pixelout<=1'b1;
25896: pixelout<=1'b1;
25897: pixelout<=1'b1;
25898: pixelout<=1'b1;
25899: pixelout<=1'b1;
25900: pixelout<=1'b1;
25901: pixelout<=1'b1;
25902: pixelout<=1'b1;
25903: pixelout<=1'b1;
25904: pixelout<=1'b1;
25905: pixelout<=1'b1;
25906: pixelout<=1'b1;
25907: pixelout<=1'b1;
25908: pixelout<=1'b1;
25909: pixelout<=1'b1;
25910: pixelout<=1'b1;
25911: pixelout<=1'b1;
25912: pixelout<=1'b1;
25913: pixelout<=1'b1;
25914: pixelout<=1'b1;
25915: pixelout<=1'b1;
25916: pixelout<=1'b1;
25917: pixelout<=1'b1;
25918: pixelout<=1'b1;
25919: pixelout<=1'b1;
25920: pixelout<=1'b1;
25921: pixelout<=1'b1;
25922: pixelout<=1'b1;
25923: pixelout<=1'b1;
25924: pixelout<=1'b1;
25925: pixelout<=1'b1;
25926: pixelout<=1'b1;
25927: pixelout<=1'b1;
25928: pixelout<=1'b1;
25929: pixelout<=1'b1;
25930: pixelout<=1'b1;
25931: pixelout<=1'b1;
25932: pixelout<=1'b1;
25933: pixelout<=1'b1;
25934: pixelout<=1'b1;
25935: pixelout<=1'b1;
25936: pixelout<=1'b1;
25937: pixelout<=1'b1;
25938: pixelout<=1'b1;
25939: pixelout<=1'b1;
25940: pixelout<=1'b1;
25941: pixelout<=1'b1;
25942: pixelout<=1'b1;
25943: pixelout<=1'b1;
25944: pixelout<=1'b1;
25945: pixelout<=1'b1;
25946: pixelout<=1'b1;
25947: pixelout<=1'b1;
25948: pixelout<=1'b1;
25949: pixelout<=1'b1;
25950: pixelout<=1'b1;
25951: pixelout<=1'b1;
25952: pixelout<=1'b1;
25953: pixelout<=1'b1;
25954: pixelout<=1'b1;
25955: pixelout<=1'b1;
25956: pixelout<=1'b1;
25957: pixelout<=1'b1;
25958: pixelout<=1'b1;
25959: pixelout<=1'b1;
25960: pixelout<=1'b1;
25961: pixelout<=1'b1;
25962: pixelout<=1'b1;
25963: pixelout<=1'b1;
25964: pixelout<=1'b1;
25965: pixelout<=1'b1;
25966: pixelout<=1'b1;
25967: pixelout<=1'b1;
25968: pixelout<=1'b1;
25969: pixelout<=1'b1;
25970: pixelout<=1'b1;
25971: pixelout<=1'b1;
25972: pixelout<=1'b1;
25973: pixelout<=1'b1;
25974: pixelout<=1'b1;
25975: pixelout<=1'b1;
25976: pixelout<=1'b1;
25977: pixelout<=1'b1;
25978: pixelout<=1'b1;
25979: pixelout<=1'b1;
25980: pixelout<=1'b1;
25981: pixelout<=1'b1;
25982: pixelout<=1'b1;
25983: pixelout<=1'b1;
25984: pixelout<=1'b1;
25985: pixelout<=1'b1;
25986: pixelout<=1'b1;
25987: pixelout<=1'b1;
25988: pixelout<=1'b1;
25989: pixelout<=1'b1;
25990: pixelout<=1'b1;
25991: pixelout<=1'b1;
25992: pixelout<=1'b1;
25993: pixelout<=1'b1;
25994: pixelout<=1'b1;
25995: pixelout<=1'b1;
25996: pixelout<=1'b1;
25997: pixelout<=1'b1;
25998: pixelout<=1'b1;
25999: pixelout<=1'b1;
26000: pixelout<=1'b1;
26001: pixelout<=1'b1;
26002: pixelout<=1'b1;
26003: pixelout<=1'b1;
26004: pixelout<=1'b1;
26005: pixelout<=1'b1;
26006: pixelout<=1'b1;
26007: pixelout<=1'b1;
26008: pixelout<=1'b1;
26009: pixelout<=1'b1;
26010: pixelout<=1'b1;
26011: pixelout<=1'b1;
26012: pixelout<=1'b1;
26013: pixelout<=1'b1;
26014: pixelout<=1'b1;
26015: pixelout<=1'b1;
26016: pixelout<=1'b0;
26017: pixelout<=1'b1;
26018: pixelout<=1'b1;
26019: pixelout<=1'b1;
26020: pixelout<=1'b1;
26021: pixelout<=1'b1;
26022: pixelout<=1'b1;
26023: pixelout<=1'b1;
26024: pixelout<=1'b1;
26025: pixelout<=1'b1;
26026: pixelout<=1'b1;
26027: pixelout<=1'b1;
26028: pixelout<=1'b1;
26029: pixelout<=1'b1;
26030: pixelout<=1'b1;
26031: pixelout<=1'b1;
26032: pixelout<=1'b1;
26033: pixelout<=1'b1;
26034: pixelout<=1'b1;
26035: pixelout<=1'b1;
26036: pixelout<=1'b1;
26037: pixelout<=1'b1;
26038: pixelout<=1'b1;
26039: pixelout<=1'b1;
26040: pixelout<=1'b1;
26041: pixelout<=1'b1;
26042: pixelout<=1'b1;
26043: pixelout<=1'b1;
26044: pixelout<=1'b1;
26045: pixelout<=1'b1;
26046: pixelout<=1'b1;
26047: pixelout<=1'b1;
26048: pixelout<=1'b1;
26049: pixelout<=1'b1;
26050: pixelout<=1'b1;
26051: pixelout<=1'b1;
26052: pixelout<=1'b1;
26053: pixelout<=1'b1;
26054: pixelout<=1'b1;
26055: pixelout<=1'b1;
26056: pixelout<=1'b1;
26057: pixelout<=1'b1;
26058: pixelout<=1'b1;
26059: pixelout<=1'b1;
26060: pixelout<=1'b1;
26061: pixelout<=1'b1;
26062: pixelout<=1'b1;
26063: pixelout<=1'b1;
26064: pixelout<=1'b1;
26065: pixelout<=1'b1;
26066: pixelout<=1'b1;
26067: pixelout<=1'b1;
26068: pixelout<=1'b1;
26069: pixelout<=1'b1;
26070: pixelout<=1'b1;
26071: pixelout<=1'b1;
26072: pixelout<=1'b1;
26073: pixelout<=1'b1;
26074: pixelout<=1'b1;
26075: pixelout<=1'b1;
26076: pixelout<=1'b1;
26077: pixelout<=1'b1;
26078: pixelout<=1'b1;
26079: pixelout<=1'b1;
26080: pixelout<=1'b1;
26081: pixelout<=1'b1;
26082: pixelout<=1'b1;
26083: pixelout<=1'b1;
26084: pixelout<=1'b1;
26085: pixelout<=1'b1;
26086: pixelout<=1'b1;
26087: pixelout<=1'b1;
26088: pixelout<=1'b1;
26089: pixelout<=1'b1;
26090: pixelout<=1'b1;
26091: pixelout<=1'b1;
26092: pixelout<=1'b1;
26093: pixelout<=1'b1;
26094: pixelout<=1'b1;
26095: pixelout<=1'b1;
26096: pixelout<=1'b1;
26097: pixelout<=1'b1;
26098: pixelout<=1'b1;
26099: pixelout<=1'b1;
26100: pixelout<=1'b1;
26101: pixelout<=1'b1;
26102: pixelout<=1'b1;
26103: pixelout<=1'b1;
26104: pixelout<=1'b1;
26105: pixelout<=1'b1;
26106: pixelout<=1'b1;
26107: pixelout<=1'b1;
26108: pixelout<=1'b1;
26109: pixelout<=1'b1;
26110: pixelout<=1'b1;
26111: pixelout<=1'b1;
26112: pixelout<=1'b1;
26113: pixelout<=1'b1;
26114: pixelout<=1'b1;
26115: pixelout<=1'b1;
26116: pixelout<=1'b1;
26117: pixelout<=1'b1;
26118: pixelout<=1'b1;
26119: pixelout<=1'b1;
26120: pixelout<=1'b1;
26121: pixelout<=1'b1;
26122: pixelout<=1'b1;
26123: pixelout<=1'b1;
26124: pixelout<=1'b1;
26125: pixelout<=1'b1;
26126: pixelout<=1'b1;
26127: pixelout<=1'b1;
26128: pixelout<=1'b1;
26129: pixelout<=1'b1;
26130: pixelout<=1'b1;
26131: pixelout<=1'b1;
26132: pixelout<=1'b1;
26133: pixelout<=1'b1;
26134: pixelout<=1'b1;
26135: pixelout<=1'b1;
26136: pixelout<=1'b1;
26137: pixelout<=1'b1;
26138: pixelout<=1'b1;
26139: pixelout<=1'b1;
26140: pixelout<=1'b1;
26141: pixelout<=1'b1;
26142: pixelout<=1'b1;
26143: pixelout<=1'b1;
26144: pixelout<=1'b1;
26145: pixelout<=1'b1;
26146: pixelout<=1'b1;
26147: pixelout<=1'b1;
26148: pixelout<=1'b1;
26149: pixelout<=1'b1;
26150: pixelout<=1'b1;
26151: pixelout<=1'b1;
26152: pixelout<=1'b1;
26153: pixelout<=1'b1;
26154: pixelout<=1'b1;
26155: pixelout<=1'b1;
26156: pixelout<=1'b1;
26157: pixelout<=1'b1;
26158: pixelout<=1'b1;
26159: pixelout<=1'b1;
26160: pixelout<=1'b1;
26161: pixelout<=1'b1;
26162: pixelout<=1'b1;
26163: pixelout<=1'b1;
26164: pixelout<=1'b1;
26165: pixelout<=1'b1;
26166: pixelout<=1'b1;
26167: pixelout<=1'b1;
26168: pixelout<=1'b1;
26169: pixelout<=1'b1;
26170: pixelout<=1'b1;
26171: pixelout<=1'b1;
26172: pixelout<=1'b1;
26173: pixelout<=1'b1;
26174: pixelout<=1'b1;
26175: pixelout<=1'b1;
26176: pixelout<=1'b1;
26177: pixelout<=1'b1;
26178: pixelout<=1'b1;
26179: pixelout<=1'b1;
26180: pixelout<=1'b1;
26181: pixelout<=1'b1;
26182: pixelout<=1'b1;
26183: pixelout<=1'b1;
26184: pixelout<=1'b1;
26185: pixelout<=1'b1;
26186: pixelout<=1'b1;
26187: pixelout<=1'b1;
26188: pixelout<=1'b1;
26189: pixelout<=1'b1;
26190: pixelout<=1'b1;
26191: pixelout<=1'b1;
26192: pixelout<=1'b1;
26193: pixelout<=1'b1;
26194: pixelout<=1'b1;
26195: pixelout<=1'b1;
26196: pixelout<=1'b1;
26197: pixelout<=1'b1;
26198: pixelout<=1'b1;
26199: pixelout<=1'b1;
26200: pixelout<=1'b1;
26201: pixelout<=1'b1;
26202: pixelout<=1'b1;
26203: pixelout<=1'b1;
26204: pixelout<=1'b1;
26205: pixelout<=1'b1;
26206: pixelout<=1'b1;
26207: pixelout<=1'b1;
26208: pixelout<=1'b1;
26209: pixelout<=1'b1;
26210: pixelout<=1'b1;
26211: pixelout<=1'b1;
26212: pixelout<=1'b1;
26213: pixelout<=1'b1;
26214: pixelout<=1'b1;
26215: pixelout<=1'b1;
26216: pixelout<=1'b1;
26217: pixelout<=1'b1;
26218: pixelout<=1'b1;
26219: pixelout<=1'b1;
26220: pixelout<=1'b1;
26221: pixelout<=1'b1;
26222: pixelout<=1'b1;
26223: pixelout<=1'b1;
26224: pixelout<=1'b1;
26225: pixelout<=1'b1;
26226: pixelout<=1'b1;
26227: pixelout<=1'b1;
26228: pixelout<=1'b1;
26229: pixelout<=1'b1;
26230: pixelout<=1'b1;
26231: pixelout<=1'b1;
26232: pixelout<=1'b1;
26233: pixelout<=1'b1;
26234: pixelout<=1'b1;
26235: pixelout<=1'b1;
26236: pixelout<=1'b1;
26237: pixelout<=1'b1;
26238: pixelout<=1'b1;
26239: pixelout<=1'b1;
26240: pixelout<=1'b1;
26241: pixelout<=1'b1;
26242: pixelout<=1'b1;
26243: pixelout<=1'b1;
26244: pixelout<=1'b1;
26245: pixelout<=1'b1;
26246: pixelout<=1'b1;
26247: pixelout<=1'b1;
26248: pixelout<=1'b1;
26249: pixelout<=1'b1;
26250: pixelout<=1'b1;
26251: pixelout<=1'b1;
26252: pixelout<=1'b1;
26253: pixelout<=1'b1;
26254: pixelout<=1'b1;
26255: pixelout<=1'b0;
26256: pixelout<=1'b1;
26257: pixelout<=1'b1;
26258: pixelout<=1'b1;
26259: pixelout<=1'b1;
26260: pixelout<=1'b1;
26261: pixelout<=1'b1;
26262: pixelout<=1'b1;
26263: pixelout<=1'b1;
26264: pixelout<=1'b1;
26265: pixelout<=1'b1;
26266: pixelout<=1'b1;
26267: pixelout<=1'b1;
26268: pixelout<=1'b1;
26269: pixelout<=1'b1;
26270: pixelout<=1'b1;
26271: pixelout<=1'b1;
26272: pixelout<=1'b1;
26273: pixelout<=1'b1;
26274: pixelout<=1'b1;
26275: pixelout<=1'b1;
26276: pixelout<=1'b1;
26277: pixelout<=1'b1;
26278: pixelout<=1'b1;
26279: pixelout<=1'b1;
26280: pixelout<=1'b1;
26281: pixelout<=1'b1;
26282: pixelout<=1'b1;
26283: pixelout<=1'b1;
26284: pixelout<=1'b1;
26285: pixelout<=1'b1;
26286: pixelout<=1'b1;
26287: pixelout<=1'b1;
26288: pixelout<=1'b1;
26289: pixelout<=1'b1;
26290: pixelout<=1'b1;
26291: pixelout<=1'b1;
26292: pixelout<=1'b1;
26293: pixelout<=1'b1;
26294: pixelout<=1'b1;
26295: pixelout<=1'b1;
26296: pixelout<=1'b1;
26297: pixelout<=1'b1;
26298: pixelout<=1'b1;
26299: pixelout<=1'b1;
26300: pixelout<=1'b1;
26301: pixelout<=1'b1;
26302: pixelout<=1'b1;
26303: pixelout<=1'b1;
26304: pixelout<=1'b1;
26305: pixelout<=1'b1;
26306: pixelout<=1'b1;
26307: pixelout<=1'b1;
26308: pixelout<=1'b1;
26309: pixelout<=1'b1;
26310: pixelout<=1'b1;
26311: pixelout<=1'b1;
26312: pixelout<=1'b1;
26313: pixelout<=1'b1;
26314: pixelout<=1'b1;
26315: pixelout<=1'b1;
26316: pixelout<=1'b1;
26317: pixelout<=1'b1;
26318: pixelout<=1'b1;
26319: pixelout<=1'b1;
26320: pixelout<=1'b1;
26321: pixelout<=1'b1;
26322: pixelout<=1'b1;
26323: pixelout<=1'b1;
26324: pixelout<=1'b1;
26325: pixelout<=1'b1;
26326: pixelout<=1'b1;
26327: pixelout<=1'b1;
26328: pixelout<=1'b1;
26329: pixelout<=1'b1;
26330: pixelout<=1'b1;
26331: pixelout<=1'b1;
26332: pixelout<=1'b1;
26333: pixelout<=1'b1;
26334: pixelout<=1'b1;
26335: pixelout<=1'b1;
26336: pixelout<=1'b1;
26337: pixelout<=1'b1;
26338: pixelout<=1'b1;
26339: pixelout<=1'b1;
26340: pixelout<=1'b1;
26341: pixelout<=1'b1;
26342: pixelout<=1'b1;
26343: pixelout<=1'b1;
26344: pixelout<=1'b1;
26345: pixelout<=1'b1;
26346: pixelout<=1'b1;
26347: pixelout<=1'b1;
26348: pixelout<=1'b1;
26349: pixelout<=1'b1;
26350: pixelout<=1'b1;
26351: pixelout<=1'b1;
26352: pixelout<=1'b1;
26353: pixelout<=1'b1;
26354: pixelout<=1'b1;
26355: pixelout<=1'b1;
26356: pixelout<=1'b1;
26357: pixelout<=1'b1;
26358: pixelout<=1'b1;
26359: pixelout<=1'b1;
26360: pixelout<=1'b1;
26361: pixelout<=1'b1;
26362: pixelout<=1'b1;
26363: pixelout<=1'b1;
26364: pixelout<=1'b1;
26365: pixelout<=1'b1;
26366: pixelout<=1'b1;
26367: pixelout<=1'b1;
26368: pixelout<=1'b1;
26369: pixelout<=1'b1;
26370: pixelout<=1'b1;
26371: pixelout<=1'b1;
26372: pixelout<=1'b1;
26373: pixelout<=1'b1;
26374: pixelout<=1'b1;
26375: pixelout<=1'b1;
26376: pixelout<=1'b1;
26377: pixelout<=1'b1;
26378: pixelout<=1'b1;
26379: pixelout<=1'b1;
26380: pixelout<=1'b1;
26381: pixelout<=1'b1;
26382: pixelout<=1'b1;
26383: pixelout<=1'b1;
26384: pixelout<=1'b1;
26385: pixelout<=1'b1;
26386: pixelout<=1'b1;
26387: pixelout<=1'b1;
26388: pixelout<=1'b1;
26389: pixelout<=1'b1;
26390: pixelout<=1'b1;
26391: pixelout<=1'b1;
26392: pixelout<=1'b1;
26393: pixelout<=1'b1;
26394: pixelout<=1'b1;
26395: pixelout<=1'b1;
26396: pixelout<=1'b1;
26397: pixelout<=1'b1;
26398: pixelout<=1'b1;
26399: pixelout<=1'b1;
26400: pixelout<=1'b1;
26401: pixelout<=1'b1;
26402: pixelout<=1'b1;
26403: pixelout<=1'b1;
26404: pixelout<=1'b1;
26405: pixelout<=1'b1;
26406: pixelout<=1'b1;
26407: pixelout<=1'b1;
26408: pixelout<=1'b1;
26409: pixelout<=1'b1;
26410: pixelout<=1'b1;
26411: pixelout<=1'b1;
26412: pixelout<=1'b1;
26413: pixelout<=1'b1;
26414: pixelout<=1'b1;
26415: pixelout<=1'b1;
26416: pixelout<=1'b1;
26417: pixelout<=1'b1;
26418: pixelout<=1'b1;
26419: pixelout<=1'b1;
26420: pixelout<=1'b0;
26421: pixelout<=1'b0;
26422: pixelout<=1'b0;
26423: pixelout<=1'b1;
26424: pixelout<=1'b1;
26425: pixelout<=1'b1;
26426: pixelout<=1'b1;
26427: pixelout<=1'b1;
26428: pixelout<=1'b1;
26429: pixelout<=1'b1;
26430: pixelout<=1'b1;
26431: pixelout<=1'b1;
26432: pixelout<=1'b1;
26433: pixelout<=1'b1;
26434: pixelout<=1'b1;
26435: pixelout<=1'b1;
26436: pixelout<=1'b1;
26437: pixelout<=1'b1;
26438: pixelout<=1'b1;
26439: pixelout<=1'b1;
26440: pixelout<=1'b1;
26441: pixelout<=1'b1;
26442: pixelout<=1'b1;
26443: pixelout<=1'b1;
26444: pixelout<=1'b1;
26445: pixelout<=1'b1;
26446: pixelout<=1'b1;
26447: pixelout<=1'b1;
26448: pixelout<=1'b1;
26449: pixelout<=1'b1;
26450: pixelout<=1'b1;
26451: pixelout<=1'b1;
26452: pixelout<=1'b1;
26453: pixelout<=1'b1;
26454: pixelout<=1'b1;
26455: pixelout<=1'b1;
26456: pixelout<=1'b1;
26457: pixelout<=1'b1;
26458: pixelout<=1'b1;
26459: pixelout<=1'b1;
26460: pixelout<=1'b1;
26461: pixelout<=1'b1;
26462: pixelout<=1'b1;
26463: pixelout<=1'b1;
26464: pixelout<=1'b1;
26465: pixelout<=1'b1;
26466: pixelout<=1'b1;
26467: pixelout<=1'b0;
26468: pixelout<=1'b1;
26469: pixelout<=1'b1;
26470: pixelout<=1'b1;
26471: pixelout<=1'b0;
26472: pixelout<=1'b0;
26473: pixelout<=1'b1;
26474: pixelout<=1'b1;
26475: pixelout<=1'b1;
26476: pixelout<=1'b1;
26477: pixelout<=1'b1;
26478: pixelout<=1'b1;
26479: pixelout<=1'b1;
26480: pixelout<=1'b1;
26481: pixelout<=1'b1;
26482: pixelout<=1'b1;
26483: pixelout<=1'b1;
26484: pixelout<=1'b1;
26485: pixelout<=1'b1;
26486: pixelout<=1'b1;
26487: pixelout<=1'b1;
26488: pixelout<=1'b1;
26489: pixelout<=1'b1;
26490: pixelout<=1'b1;
26491: pixelout<=1'b1;
26492: pixelout<=1'b1;
26493: pixelout<=1'b1;
26494: pixelout<=1'b1;
26495: pixelout<=1'b1;
26496: pixelout<=1'b1;
26497: pixelout<=1'b1;
26498: pixelout<=1'b1;
26499: pixelout<=1'b1;
26500: pixelout<=1'b1;
26501: pixelout<=1'b1;
26502: pixelout<=1'b1;
26503: pixelout<=1'b1;
26504: pixelout<=1'b1;
26505: pixelout<=1'b1;
26506: pixelout<=1'b1;
26507: pixelout<=1'b1;
26508: pixelout<=1'b1;
26509: pixelout<=1'b1;
26510: pixelout<=1'b1;
26511: pixelout<=1'b1;
26512: pixelout<=1'b1;
26513: pixelout<=1'b1;
26514: pixelout<=1'b1;
26515: pixelout<=1'b1;
26516: pixelout<=1'b1;
26517: pixelout<=1'b1;
26518: pixelout<=1'b1;
26519: pixelout<=1'b1;
26520: pixelout<=1'b1;
26521: pixelout<=1'b1;
26522: pixelout<=1'b1;
26523: pixelout<=1'b1;
26524: pixelout<=1'b1;
26525: pixelout<=1'b1;
26526: pixelout<=1'b1;
26527: pixelout<=1'b1;
26528: pixelout<=1'b1;
26529: pixelout<=1'b1;
26530: pixelout<=1'b1;
26531: pixelout<=1'b1;
26532: pixelout<=1'b1;
26533: pixelout<=1'b1;
26534: pixelout<=1'b0;
26535: pixelout<=1'b1;
26536: pixelout<=1'b1;
26537: pixelout<=1'b1;
26538: pixelout<=1'b1;
26539: pixelout<=1'b1;
26540: pixelout<=1'b1;
26541: pixelout<=1'b1;
26542: pixelout<=1'b1;
26543: pixelout<=1'b1;
26544: pixelout<=1'b1;
26545: pixelout<=1'b1;
26546: pixelout<=1'b1;
26547: pixelout<=1'b1;
26548: pixelout<=1'b1;
26549: pixelout<=1'b1;
26550: pixelout<=1'b1;
26551: pixelout<=1'b1;
26552: pixelout<=1'b1;
26553: pixelout<=1'b1;
26554: pixelout<=1'b1;
26555: pixelout<=1'b1;
26556: pixelout<=1'b1;
26557: pixelout<=1'b1;
26558: pixelout<=1'b1;
26559: pixelout<=1'b1;
26560: pixelout<=1'b1;
26561: pixelout<=1'b1;
26562: pixelout<=1'b1;
26563: pixelout<=1'b1;
26564: pixelout<=1'b1;
26565: pixelout<=1'b1;
26566: pixelout<=1'b1;
26567: pixelout<=1'b1;
26568: pixelout<=1'b1;
26569: pixelout<=1'b1;
26570: pixelout<=1'b1;
26571: pixelout<=1'b1;
26572: pixelout<=1'b1;
26573: pixelout<=1'b1;
26574: pixelout<=1'b1;
26575: pixelout<=1'b1;
26576: pixelout<=1'b1;
26577: pixelout<=1'b1;
26578: pixelout<=1'b1;
26579: pixelout<=1'b1;
26580: pixelout<=1'b1;
26581: pixelout<=1'b1;
26582: pixelout<=1'b1;
26583: pixelout<=1'b1;
26584: pixelout<=1'b1;
26585: pixelout<=1'b1;
26586: pixelout<=1'b1;
26587: pixelout<=1'b1;
26588: pixelout<=1'b1;
26589: pixelout<=1'b1;
26590: pixelout<=1'b0;
26591: pixelout<=1'b1;
26592: pixelout<=1'b1;
26593: pixelout<=1'b1;
26594: pixelout<=1'b0;
26595: pixelout<=1'b1;
26596: pixelout<=1'b1;
26597: pixelout<=1'b1;
26598: pixelout<=1'b1;
26599: pixelout<=1'b1;
26600: pixelout<=1'b1;
26601: pixelout<=1'b1;
26602: pixelout<=1'b1;
26603: pixelout<=1'b1;
26604: pixelout<=1'b1;
26605: pixelout<=1'b1;
26606: pixelout<=1'b1;
26607: pixelout<=1'b1;
26608: pixelout<=1'b1;
26609: pixelout<=1'b1;
26610: pixelout<=1'b1;
26611: pixelout<=1'b1;
26612: pixelout<=1'b1;
26613: pixelout<=1'b1;
26614: pixelout<=1'b1;
26615: pixelout<=1'b1;
26616: pixelout<=1'b1;
26617: pixelout<=1'b1;
26618: pixelout<=1'b1;
26619: pixelout<=1'b1;
26620: pixelout<=1'b1;
26621: pixelout<=1'b1;
26622: pixelout<=1'b1;
26623: pixelout<=1'b1;
26624: pixelout<=1'b1;
26625: pixelout<=1'b1;
26626: pixelout<=1'b1;
26627: pixelout<=1'b1;
26628: pixelout<=1'b1;
26629: pixelout<=1'b1;
26630: pixelout<=1'b1;
26631: pixelout<=1'b1;
26632: pixelout<=1'b1;
26633: pixelout<=1'b1;
26634: pixelout<=1'b1;
26635: pixelout<=1'b1;
26636: pixelout<=1'b1;
26637: pixelout<=1'b1;
26638: pixelout<=1'b1;
26639: pixelout<=1'b1;
26640: pixelout<=1'b1;
26641: pixelout<=1'b1;
26642: pixelout<=1'b1;
26643: pixelout<=1'b1;
26644: pixelout<=1'b1;
26645: pixelout<=1'b1;
26646: pixelout<=1'b1;
26647: pixelout<=1'b1;
26648: pixelout<=1'b1;
26649: pixelout<=1'b1;
26650: pixelout<=1'b1;
26651: pixelout<=1'b1;
26652: pixelout<=1'b1;
26653: pixelout<=1'b1;
26654: pixelout<=1'b1;
26655: pixelout<=1'b1;
26656: pixelout<=1'b1;
26657: pixelout<=1'b1;
26658: pixelout<=1'b1;
26659: pixelout<=1'b0;
26660: pixelout<=1'b1;
26661: pixelout<=1'b1;
26662: pixelout<=1'b1;
26663: pixelout<=1'b1;
26664: pixelout<=1'b1;
26665: pixelout<=1'b1;
26666: pixelout<=1'b1;
26667: pixelout<=1'b1;
26668: pixelout<=1'b1;
26669: pixelout<=1'b1;
26670: pixelout<=1'b1;
26671: pixelout<=1'b1;
26672: pixelout<=1'b1;
26673: pixelout<=1'b1;
26674: pixelout<=1'b1;
26675: pixelout<=1'b1;
26676: pixelout<=1'b1;
26677: pixelout<=1'b1;
26678: pixelout<=1'b1;
26679: pixelout<=1'b1;
26680: pixelout<=1'b1;
26681: pixelout<=1'b1;
26682: pixelout<=1'b1;
26683: pixelout<=1'b1;
26684: pixelout<=1'b1;
26685: pixelout<=1'b1;
26686: pixelout<=1'b1;
26687: pixelout<=1'b1;
26688: pixelout<=1'b1;
26689: pixelout<=1'b1;
26690: pixelout<=1'b1;
26691: pixelout<=1'b1;
26692: pixelout<=1'b1;
26693: pixelout<=1'b1;
26694: pixelout<=1'b1;
26695: pixelout<=1'b1;
26696: pixelout<=1'b1;
26697: pixelout<=1'b1;
26698: pixelout<=1'b1;
26699: pixelout<=1'b1;
26700: pixelout<=1'b1;
26701: pixelout<=1'b1;
26702: pixelout<=1'b1;
26703: pixelout<=1'b1;
26704: pixelout<=1'b1;
26705: pixelout<=1'b1;
26706: pixelout<=1'b1;
26707: pixelout<=1'b1;
26708: pixelout<=1'b1;
26709: pixelout<=1'b1;
26710: pixelout<=1'b0;
26711: pixelout<=1'b1;
26712: pixelout<=1'b1;
26713: pixelout<=1'b1;
26714: pixelout<=1'b1;
26715: pixelout<=1'b1;
26716: pixelout<=1'b1;
26717: pixelout<=1'b1;
26718: pixelout<=1'b1;
26719: pixelout<=1'b1;
26720: pixelout<=1'b1;
26721: pixelout<=1'b1;
26722: pixelout<=1'b1;
26723: pixelout<=1'b1;
26724: pixelout<=1'b1;
26725: pixelout<=1'b1;
26726: pixelout<=1'b1;
26727: pixelout<=1'b1;
26728: pixelout<=1'b1;
26729: pixelout<=1'b1;
26730: pixelout<=1'b1;
26731: pixelout<=1'b1;
26732: pixelout<=1'b1;
26733: pixelout<=1'b1;
26734: pixelout<=1'b1;
26735: pixelout<=1'b1;
26736: pixelout<=1'b1;
26737: pixelout<=1'b1;
26738: pixelout<=1'b1;
26739: pixelout<=1'b1;
26740: pixelout<=1'b1;
26741: pixelout<=1'b1;
26742: pixelout<=1'b1;
26743: pixelout<=1'b1;
26744: pixelout<=1'b1;
26745: pixelout<=1'b1;
26746: pixelout<=1'b1;
26747: pixelout<=1'b1;
26748: pixelout<=1'b1;
26749: pixelout<=1'b1;
26750: pixelout<=1'b1;
26751: pixelout<=1'b1;
26752: pixelout<=1'b1;
26753: pixelout<=1'b1;
26754: pixelout<=1'b1;
26755: pixelout<=1'b1;
26756: pixelout<=1'b1;
26757: pixelout<=1'b1;
26758: pixelout<=1'b1;
26759: pixelout<=1'b1;
26760: pixelout<=1'b1;
26761: pixelout<=1'b1;
26762: pixelout<=1'b1;
26763: pixelout<=1'b1;
26764: pixelout<=1'b1;
26765: pixelout<=1'b1;
26766: pixelout<=1'b1;
26767: pixelout<=1'b1;
26768: pixelout<=1'b1;
26769: pixelout<=1'b1;
26770: pixelout<=1'b1;
26771: pixelout<=1'b1;
26772: pixelout<=1'b1;
26773: pixelout<=1'b1;
26774: pixelout<=1'b0;
26775: pixelout<=1'b1;
26776: pixelout<=1'b1;
26777: pixelout<=1'b1;
26778: pixelout<=1'b1;
26779: pixelout<=1'b1;
26780: pixelout<=1'b1;
26781: pixelout<=1'b1;
26782: pixelout<=1'b1;
26783: pixelout<=1'b1;
26784: pixelout<=1'b1;
26785: pixelout<=1'b1;
26786: pixelout<=1'b1;
26787: pixelout<=1'b1;
26788: pixelout<=1'b1;
26789: pixelout<=1'b0;
26790: pixelout<=1'b1;
26791: pixelout<=1'b1;
26792: pixelout<=1'b1;
26793: pixelout<=1'b1;
26794: pixelout<=1'b1;
26795: pixelout<=1'b1;
26796: pixelout<=1'b1;
26797: pixelout<=1'b1;
26798: pixelout<=1'b1;
26799: pixelout<=1'b1;
26800: pixelout<=1'b1;
26801: pixelout<=1'b1;
26802: pixelout<=1'b1;
26803: pixelout<=1'b1;
26804: pixelout<=1'b1;
26805: pixelout<=1'b1;
26806: pixelout<=1'b1;
26807: pixelout<=1'b1;
26808: pixelout<=1'b1;
26809: pixelout<=1'b1;
26810: pixelout<=1'b1;
26811: pixelout<=1'b1;
26812: pixelout<=1'b1;
26813: pixelout<=1'b1;
26814: pixelout<=1'b1;
26815: pixelout<=1'b1;
26816: pixelout<=1'b1;
26817: pixelout<=1'b1;
26818: pixelout<=1'b1;
26819: pixelout<=1'b1;
26820: pixelout<=1'b1;
26821: pixelout<=1'b1;
26822: pixelout<=1'b1;
26823: pixelout<=1'b1;
26824: pixelout<=1'b1;
26825: pixelout<=1'b1;
26826: pixelout<=1'b1;
26827: pixelout<=1'b1;
26828: pixelout<=1'b1;
26829: pixelout<=1'b1;
26830: pixelout<=1'b0;
26831: pixelout<=1'b1;
26832: pixelout<=1'b1;
26833: pixelout<=1'b1;
26834: pixelout<=1'b0;
26835: pixelout<=1'b1;
26836: pixelout<=1'b1;
26837: pixelout<=1'b1;
26838: pixelout<=1'b1;
26839: pixelout<=1'b1;
26840: pixelout<=1'b1;
26841: pixelout<=1'b1;
26842: pixelout<=1'b1;
26843: pixelout<=1'b1;
26844: pixelout<=1'b1;
26845: pixelout<=1'b1;
26846: pixelout<=1'b1;
26847: pixelout<=1'b1;
26848: pixelout<=1'b1;
26849: pixelout<=1'b1;
26850: pixelout<=1'b1;
26851: pixelout<=1'b1;
26852: pixelout<=1'b1;
26853: pixelout<=1'b1;
26854: pixelout<=1'b1;
26855: pixelout<=1'b1;
26856: pixelout<=1'b1;
26857: pixelout<=1'b1;
26858: pixelout<=1'b1;
26859: pixelout<=1'b1;
26860: pixelout<=1'b1;
26861: pixelout<=1'b1;
26862: pixelout<=1'b1;
26863: pixelout<=1'b1;
26864: pixelout<=1'b1;
26865: pixelout<=1'b1;
26866: pixelout<=1'b1;
26867: pixelout<=1'b1;
26868: pixelout<=1'b1;
26869: pixelout<=1'b1;
26870: pixelout<=1'b1;
26871: pixelout<=1'b1;
26872: pixelout<=1'b1;
26873: pixelout<=1'b1;
26874: pixelout<=1'b1;
26875: pixelout<=1'b1;
26876: pixelout<=1'b1;
26877: pixelout<=1'b1;
26878: pixelout<=1'b1;
26879: pixelout<=1'b1;
26880: pixelout<=1'b1;
26881: pixelout<=1'b1;
26882: pixelout<=1'b1;
26883: pixelout<=1'b1;
26884: pixelout<=1'b1;
26885: pixelout<=1'b1;
26886: pixelout<=1'b1;
26887: pixelout<=1'b1;
26888: pixelout<=1'b1;
26889: pixelout<=1'b1;
26890: pixelout<=1'b1;
26891: pixelout<=1'b1;
26892: pixelout<=1'b1;
26893: pixelout<=1'b1;
26894: pixelout<=1'b1;
26895: pixelout<=1'b1;
26896: pixelout<=1'b1;
26897: pixelout<=1'b1;
26898: pixelout<=1'b1;
26899: pixelout<=1'b0;
26900: pixelout<=1'b1;
26901: pixelout<=1'b1;
26902: pixelout<=1'b1;
26903: pixelout<=1'b1;
26904: pixelout<=1'b1;
26905: pixelout<=1'b1;
26906: pixelout<=1'b1;
26907: pixelout<=1'b1;
26908: pixelout<=1'b1;
26909: pixelout<=1'b1;
26910: pixelout<=1'b1;
26911: pixelout<=1'b1;
26912: pixelout<=1'b1;
26913: pixelout<=1'b1;
26914: pixelout<=1'b1;
26915: pixelout<=1'b1;
26916: pixelout<=1'b1;
26917: pixelout<=1'b1;
26918: pixelout<=1'b1;
26919: pixelout<=1'b1;
26920: pixelout<=1'b1;
26921: pixelout<=1'b1;
26922: pixelout<=1'b1;
26923: pixelout<=1'b1;
26924: pixelout<=1'b1;
26925: pixelout<=1'b1;
26926: pixelout<=1'b1;
26927: pixelout<=1'b1;
26928: pixelout<=1'b1;
26929: pixelout<=1'b1;
26930: pixelout<=1'b1;
26931: pixelout<=1'b1;
26932: pixelout<=1'b1;
26933: pixelout<=1'b1;
26934: pixelout<=1'b1;
26935: pixelout<=1'b1;
26936: pixelout<=1'b1;
26937: pixelout<=1'b1;
26938: pixelout<=1'b1;
26939: pixelout<=1'b1;
26940: pixelout<=1'b1;
26941: pixelout<=1'b1;
26942: pixelout<=1'b1;
26943: pixelout<=1'b1;
26944: pixelout<=1'b1;
26945: pixelout<=1'b1;
26946: pixelout<=1'b1;
26947: pixelout<=1'b1;
26948: pixelout<=1'b1;
26949: pixelout<=1'b1;
26950: pixelout<=1'b0;
26951: pixelout<=1'b1;
26952: pixelout<=1'b1;
26953: pixelout<=1'b1;
26954: pixelout<=1'b1;
26955: pixelout<=1'b1;
26956: pixelout<=1'b1;
26957: pixelout<=1'b1;
26958: pixelout<=1'b1;
26959: pixelout<=1'b1;
26960: pixelout<=1'b1;
26961: pixelout<=1'b1;
26962: pixelout<=1'b1;
26963: pixelout<=1'b1;
26964: pixelout<=1'b1;
26965: pixelout<=1'b1;
26966: pixelout<=1'b1;
26967: pixelout<=1'b1;
26968: pixelout<=1'b1;
26969: pixelout<=1'b1;
26970: pixelout<=1'b1;
26971: pixelout<=1'b1;
26972: pixelout<=1'b1;
26973: pixelout<=1'b1;
26974: pixelout<=1'b1;
26975: pixelout<=1'b1;
26976: pixelout<=1'b1;
26977: pixelout<=1'b1;
26978: pixelout<=1'b1;
26979: pixelout<=1'b1;
26980: pixelout<=1'b1;
26981: pixelout<=1'b1;
26982: pixelout<=1'b1;
26983: pixelout<=1'b1;
26984: pixelout<=1'b1;
26985: pixelout<=1'b1;
26986: pixelout<=1'b1;
26987: pixelout<=1'b1;
26988: pixelout<=1'b1;
26989: pixelout<=1'b1;
26990: pixelout<=1'b1;
26991: pixelout<=1'b1;
26992: pixelout<=1'b1;
26993: pixelout<=1'b1;
26994: pixelout<=1'b1;
26995: pixelout<=1'b1;
26996: pixelout<=1'b1;
26997: pixelout<=1'b1;
26998: pixelout<=1'b1;
26999: pixelout<=1'b1;
27000: pixelout<=1'b1;
27001: pixelout<=1'b1;
27002: pixelout<=1'b1;
27003: pixelout<=1'b1;
27004: pixelout<=1'b1;
27005: pixelout<=1'b1;
27006: pixelout<=1'b1;
27007: pixelout<=1'b1;
27008: pixelout<=1'b1;
27009: pixelout<=1'b1;
27010: pixelout<=1'b1;
27011: pixelout<=1'b1;
27012: pixelout<=1'b1;
27013: pixelout<=1'b1;
27014: pixelout<=1'b0;
27015: pixelout<=1'b1;
27016: pixelout<=1'b1;
27017: pixelout<=1'b1;
27018: pixelout<=1'b1;
27019: pixelout<=1'b1;
27020: pixelout<=1'b1;
27021: pixelout<=1'b1;
27022: pixelout<=1'b1;
27023: pixelout<=1'b1;
27024: pixelout<=1'b1;
27025: pixelout<=1'b1;
27026: pixelout<=1'b1;
27027: pixelout<=1'b1;
27028: pixelout<=1'b1;
27029: pixelout<=1'b0;
27030: pixelout<=1'b1;
27031: pixelout<=1'b1;
27032: pixelout<=1'b1;
27033: pixelout<=1'b1;
27034: pixelout<=1'b1;
27035: pixelout<=1'b1;
27036: pixelout<=1'b1;
27037: pixelout<=1'b1;
27038: pixelout<=1'b1;
27039: pixelout<=1'b1;
27040: pixelout<=1'b1;
27041: pixelout<=1'b1;
27042: pixelout<=1'b1;
27043: pixelout<=1'b1;
27044: pixelout<=1'b1;
27045: pixelout<=1'b1;
27046: pixelout<=1'b1;
27047: pixelout<=1'b1;
27048: pixelout<=1'b1;
27049: pixelout<=1'b1;
27050: pixelout<=1'b1;
27051: pixelout<=1'b1;
27052: pixelout<=1'b1;
27053: pixelout<=1'b1;
27054: pixelout<=1'b1;
27055: pixelout<=1'b1;
27056: pixelout<=1'b1;
27057: pixelout<=1'b1;
27058: pixelout<=1'b1;
27059: pixelout<=1'b1;
27060: pixelout<=1'b1;
27061: pixelout<=1'b1;
27062: pixelout<=1'b1;
27063: pixelout<=1'b1;
27064: pixelout<=1'b1;
27065: pixelout<=1'b1;
27066: pixelout<=1'b1;
27067: pixelout<=1'b1;
27068: pixelout<=1'b1;
27069: pixelout<=1'b1;
27070: pixelout<=1'b0;
27071: pixelout<=1'b1;
27072: pixelout<=1'b1;
27073: pixelout<=1'b1;
27074: pixelout<=1'b0;
27075: pixelout<=1'b1;
27076: pixelout<=1'b1;
27077: pixelout<=1'b1;
27078: pixelout<=1'b1;
27079: pixelout<=1'b1;
27080: pixelout<=1'b1;
27081: pixelout<=1'b1;
27082: pixelout<=1'b1;
27083: pixelout<=1'b1;
27084: pixelout<=1'b1;
27085: pixelout<=1'b1;
27086: pixelout<=1'b1;
27087: pixelout<=1'b1;
27088: pixelout<=1'b1;
27089: pixelout<=1'b1;
27090: pixelout<=1'b1;
27091: pixelout<=1'b1;
27092: pixelout<=1'b1;
27093: pixelout<=1'b1;
27094: pixelout<=1'b1;
27095: pixelout<=1'b1;
27096: pixelout<=1'b1;
27097: pixelout<=1'b1;
27098: pixelout<=1'b1;
27099: pixelout<=1'b1;
27100: pixelout<=1'b1;
27101: pixelout<=1'b1;
27102: pixelout<=1'b1;
27103: pixelout<=1'b1;
27104: pixelout<=1'b1;
27105: pixelout<=1'b1;
27106: pixelout<=1'b1;
27107: pixelout<=1'b1;
27108: pixelout<=1'b1;
27109: pixelout<=1'b1;
27110: pixelout<=1'b1;
27111: pixelout<=1'b1;
27112: pixelout<=1'b1;
27113: pixelout<=1'b1;
27114: pixelout<=1'b1;
27115: pixelout<=1'b1;
27116: pixelout<=1'b1;
27117: pixelout<=1'b1;
27118: pixelout<=1'b1;
27119: pixelout<=1'b1;
27120: pixelout<=1'b1;
27121: pixelout<=1'b1;
27122: pixelout<=1'b1;
27123: pixelout<=1'b1;
27124: pixelout<=1'b1;
27125: pixelout<=1'b1;
27126: pixelout<=1'b1;
27127: pixelout<=1'b1;
27128: pixelout<=1'b1;
27129: pixelout<=1'b1;
27130: pixelout<=1'b1;
27131: pixelout<=1'b1;
27132: pixelout<=1'b1;
27133: pixelout<=1'b1;
27134: pixelout<=1'b1;
27135: pixelout<=1'b1;
27136: pixelout<=1'b1;
27137: pixelout<=1'b1;
27138: pixelout<=1'b1;
27139: pixelout<=1'b0;
27140: pixelout<=1'b1;
27141: pixelout<=1'b1;
27142: pixelout<=1'b1;
27143: pixelout<=1'b1;
27144: pixelout<=1'b1;
27145: pixelout<=1'b1;
27146: pixelout<=1'b1;
27147: pixelout<=1'b0;
27148: pixelout<=1'b0;
27149: pixelout<=1'b1;
27150: pixelout<=1'b1;
27151: pixelout<=1'b1;
27152: pixelout<=1'b0;
27153: pixelout<=1'b0;
27154: pixelout<=1'b1;
27155: pixelout<=1'b1;
27156: pixelout<=1'b1;
27157: pixelout<=1'b1;
27158: pixelout<=1'b0;
27159: pixelout<=1'b0;
27160: pixelout<=1'b0;
27161: pixelout<=1'b1;
27162: pixelout<=1'b1;
27163: pixelout<=1'b0;
27164: pixelout<=1'b1;
27165: pixelout<=1'b0;
27166: pixelout<=1'b0;
27167: pixelout<=1'b1;
27168: pixelout<=1'b1;
27169: pixelout<=1'b1;
27170: pixelout<=1'b0;
27171: pixelout<=1'b0;
27172: pixelout<=1'b0;
27173: pixelout<=1'b1;
27174: pixelout<=1'b1;
27175: pixelout<=1'b0;
27176: pixelout<=1'b0;
27177: pixelout<=1'b0;
27178: pixelout<=1'b1;
27179: pixelout<=1'b1;
27180: pixelout<=1'b0;
27181: pixelout<=1'b0;
27182: pixelout<=1'b0;
27183: pixelout<=1'b0;
27184: pixelout<=1'b1;
27185: pixelout<=1'b1;
27186: pixelout<=1'b1;
27187: pixelout<=1'b0;
27188: pixelout<=1'b1;
27189: pixelout<=1'b0;
27190: pixelout<=1'b0;
27191: pixelout<=1'b0;
27192: pixelout<=1'b0;
27193: pixelout<=1'b1;
27194: pixelout<=1'b1;
27195: pixelout<=1'b1;
27196: pixelout<=1'b0;
27197: pixelout<=1'b1;
27198: pixelout<=1'b1;
27199: pixelout<=1'b1;
27200: pixelout<=1'b1;
27201: pixelout<=1'b1;
27202: pixelout<=1'b1;
27203: pixelout<=1'b1;
27204: pixelout<=1'b0;
27205: pixelout<=1'b0;
27206: pixelout<=1'b1;
27207: pixelout<=1'b1;
27208: pixelout<=1'b1;
27209: pixelout<=1'b0;
27210: pixelout<=1'b1;
27211: pixelout<=1'b1;
27212: pixelout<=1'b0;
27213: pixelout<=1'b1;
27214: pixelout<=1'b1;
27215: pixelout<=1'b1;
27216: pixelout<=1'b1;
27217: pixelout<=1'b1;
27218: pixelout<=1'b0;
27219: pixelout<=1'b1;
27220: pixelout<=1'b1;
27221: pixelout<=1'b0;
27222: pixelout<=1'b1;
27223: pixelout<=1'b1;
27224: pixelout<=1'b1;
27225: pixelout<=1'b0;
27226: pixelout<=1'b0;
27227: pixelout<=1'b1;
27228: pixelout<=1'b1;
27229: pixelout<=1'b1;
27230: pixelout<=1'b1;
27231: pixelout<=1'b1;
27232: pixelout<=1'b1;
27233: pixelout<=1'b0;
27234: pixelout<=1'b0;
27235: pixelout<=1'b0;
27236: pixelout<=1'b1;
27237: pixelout<=1'b1;
27238: pixelout<=1'b0;
27239: pixelout<=1'b1;
27240: pixelout<=1'b0;
27241: pixelout<=1'b0;
27242: pixelout<=1'b1;
27243: pixelout<=1'b1;
27244: pixelout<=1'b1;
27245: pixelout<=1'b0;
27246: pixelout<=1'b0;
27247: pixelout<=1'b0;
27248: pixelout<=1'b1;
27249: pixelout<=1'b1;
27250: pixelout<=1'b1;
27251: pixelout<=1'b0;
27252: pixelout<=1'b0;
27253: pixelout<=1'b0;
27254: pixelout<=1'b0;
27255: pixelout<=1'b1;
27256: pixelout<=1'b0;
27257: pixelout<=1'b1;
27258: pixelout<=1'b1;
27259: pixelout<=1'b0;
27260: pixelout<=1'b1;
27261: pixelout<=1'b1;
27262: pixelout<=1'b1;
27263: pixelout<=1'b0;
27264: pixelout<=1'b0;
27265: pixelout<=1'b0;
27266: pixelout<=1'b0;
27267: pixelout<=1'b1;
27268: pixelout<=1'b1;
27269: pixelout<=1'b0;
27270: pixelout<=1'b0;
27271: pixelout<=1'b0;
27272: pixelout<=1'b1;
27273: pixelout<=1'b1;
27274: pixelout<=1'b1;
27275: pixelout<=1'b1;
27276: pixelout<=1'b0;
27277: pixelout<=1'b0;
27278: pixelout<=1'b1;
27279: pixelout<=1'b1;
27280: pixelout<=1'b1;
27281: pixelout<=1'b1;
27282: pixelout<=1'b0;
27283: pixelout<=1'b0;
27284: pixelout<=1'b0;
27285: pixelout<=1'b1;
27286: pixelout<=1'b1;
27287: pixelout<=1'b1;
27288: pixelout<=1'b1;
27289: pixelout<=1'b1;
27290: pixelout<=1'b1;
27291: pixelout<=1'b1;
27292: pixelout<=1'b1;
27293: pixelout<=1'b1;
27294: pixelout<=1'b1;
27295: pixelout<=1'b1;
27296: pixelout<=1'b0;
27297: pixelout<=1'b0;
27298: pixelout<=1'b0;
27299: pixelout<=1'b1;
27300: pixelout<=1'b1;
27301: pixelout<=1'b0;
27302: pixelout<=1'b0;
27303: pixelout<=1'b1;
27304: pixelout<=1'b1;
27305: pixelout<=1'b1;
27306: pixelout<=1'b1;
27307: pixelout<=1'b0;
27308: pixelout<=1'b0;
27309: pixelout<=1'b0;
27310: pixelout<=1'b0;
27311: pixelout<=1'b1;
27312: pixelout<=1'b1;
27313: pixelout<=1'b1;
27314: pixelout<=1'b0;
27315: pixelout<=1'b0;
27316: pixelout<=1'b0;
27317: pixelout<=1'b0;
27318: pixelout<=1'b1;
27319: pixelout<=1'b1;
27320: pixelout<=1'b1;
27321: pixelout<=1'b1;
27322: pixelout<=1'b0;
27323: pixelout<=1'b0;
27324: pixelout<=1'b0;
27325: pixelout<=1'b1;
27326: pixelout<=1'b1;
27327: pixelout<=1'b1;
27328: pixelout<=1'b1;
27329: pixelout<=1'b1;
27330: pixelout<=1'b1;
27331: pixelout<=1'b0;
27332: pixelout<=1'b1;
27333: pixelout<=1'b1;
27334: pixelout<=1'b0;
27335: pixelout<=1'b0;
27336: pixelout<=1'b0;
27337: pixelout<=1'b1;
27338: pixelout<=1'b1;
27339: pixelout<=1'b1;
27340: pixelout<=1'b1;
27341: pixelout<=1'b1;
27342: pixelout<=1'b1;
27343: pixelout<=1'b1;
27344: pixelout<=1'b1;
27345: pixelout<=1'b1;
27346: pixelout<=1'b1;
27347: pixelout<=1'b1;
27348: pixelout<=1'b1;
27349: pixelout<=1'b1;
27350: pixelout<=1'b1;
27351: pixelout<=1'b1;
27352: pixelout<=1'b1;
27353: pixelout<=1'b1;
27354: pixelout<=1'b1;
27355: pixelout<=1'b1;
27356: pixelout<=1'b1;
27357: pixelout<=1'b1;
27358: pixelout<=1'b1;
27359: pixelout<=1'b1;
27360: pixelout<=1'b1;
27361: pixelout<=1'b1;
27362: pixelout<=1'b1;
27363: pixelout<=1'b1;
27364: pixelout<=1'b1;
27365: pixelout<=1'b1;
27366: pixelout<=1'b1;
27367: pixelout<=1'b1;
27368: pixelout<=1'b1;
27369: pixelout<=1'b1;
27370: pixelout<=1'b1;
27371: pixelout<=1'b1;
27372: pixelout<=1'b1;
27373: pixelout<=1'b1;
27374: pixelout<=1'b1;
27375: pixelout<=1'b1;
27376: pixelout<=1'b1;
27377: pixelout<=1'b1;
27378: pixelout<=1'b1;
27379: pixelout<=1'b0;
27380: pixelout<=1'b1;
27381: pixelout<=1'b1;
27382: pixelout<=1'b1;
27383: pixelout<=1'b1;
27384: pixelout<=1'b1;
27385: pixelout<=1'b0;
27386: pixelout<=1'b1;
27387: pixelout<=1'b1;
27388: pixelout<=1'b1;
27389: pixelout<=1'b1;
27390: pixelout<=1'b1;
27391: pixelout<=1'b1;
27392: pixelout<=1'b1;
27393: pixelout<=1'b1;
27394: pixelout<=1'b1;
27395: pixelout<=1'b0;
27396: pixelout<=1'b1;
27397: pixelout<=1'b0;
27398: pixelout<=1'b1;
27399: pixelout<=1'b1;
27400: pixelout<=1'b1;
27401: pixelout<=1'b0;
27402: pixelout<=1'b1;
27403: pixelout<=1'b0;
27404: pixelout<=1'b0;
27405: pixelout<=1'b1;
27406: pixelout<=1'b1;
27407: pixelout<=1'b1;
27408: pixelout<=1'b0;
27409: pixelout<=1'b1;
27410: pixelout<=1'b1;
27411: pixelout<=1'b1;
27412: pixelout<=1'b1;
27413: pixelout<=1'b1;
27414: pixelout<=1'b1;
27415: pixelout<=1'b1;
27416: pixelout<=1'b1;
27417: pixelout<=1'b1;
27418: pixelout<=1'b1;
27419: pixelout<=1'b1;
27420: pixelout<=1'b0;
27421: pixelout<=1'b1;
27422: pixelout<=1'b1;
27423: pixelout<=1'b1;
27424: pixelout<=1'b1;
27425: pixelout<=1'b1;
27426: pixelout<=1'b1;
27427: pixelout<=1'b0;
27428: pixelout<=1'b1;
27429: pixelout<=1'b1;
27430: pixelout<=1'b0;
27431: pixelout<=1'b1;
27432: pixelout<=1'b1;
27433: pixelout<=1'b1;
27434: pixelout<=1'b1;
27435: pixelout<=1'b1;
27436: pixelout<=1'b0;
27437: pixelout<=1'b1;
27438: pixelout<=1'b1;
27439: pixelout<=1'b1;
27440: pixelout<=1'b1;
27441: pixelout<=1'b1;
27442: pixelout<=1'b1;
27443: pixelout<=1'b1;
27444: pixelout<=1'b1;
27445: pixelout<=1'b1;
27446: pixelout<=1'b1;
27447: pixelout<=1'b0;
27448: pixelout<=1'b1;
27449: pixelout<=1'b0;
27450: pixelout<=1'b1;
27451: pixelout<=1'b1;
27452: pixelout<=1'b0;
27453: pixelout<=1'b1;
27454: pixelout<=1'b1;
27455: pixelout<=1'b1;
27456: pixelout<=1'b1;
27457: pixelout<=1'b1;
27458: pixelout<=1'b0;
27459: pixelout<=1'b0;
27460: pixelout<=1'b1;
27461: pixelout<=1'b1;
27462: pixelout<=1'b1;
27463: pixelout<=1'b1;
27464: pixelout<=1'b1;
27465: pixelout<=1'b1;
27466: pixelout<=1'b1;
27467: pixelout<=1'b1;
27468: pixelout<=1'b0;
27469: pixelout<=1'b1;
27470: pixelout<=1'b1;
27471: pixelout<=1'b1;
27472: pixelout<=1'b0;
27473: pixelout<=1'b1;
27474: pixelout<=1'b1;
27475: pixelout<=1'b1;
27476: pixelout<=1'b0;
27477: pixelout<=1'b1;
27478: pixelout<=1'b0;
27479: pixelout<=1'b0;
27480: pixelout<=1'b1;
27481: pixelout<=1'b1;
27482: pixelout<=1'b1;
27483: pixelout<=1'b0;
27484: pixelout<=1'b1;
27485: pixelout<=1'b1;
27486: pixelout<=1'b1;
27487: pixelout<=1'b1;
27488: pixelout<=1'b1;
27489: pixelout<=1'b1;
27490: pixelout<=1'b1;
27491: pixelout<=1'b1;
27492: pixelout<=1'b1;
27493: pixelout<=1'b1;
27494: pixelout<=1'b0;
27495: pixelout<=1'b1;
27496: pixelout<=1'b0;
27497: pixelout<=1'b1;
27498: pixelout<=1'b1;
27499: pixelout<=1'b0;
27500: pixelout<=1'b1;
27501: pixelout<=1'b1;
27502: pixelout<=1'b0;
27503: pixelout<=1'b1;
27504: pixelout<=1'b1;
27505: pixelout<=1'b1;
27506: pixelout<=1'b0;
27507: pixelout<=1'b1;
27508: pixelout<=1'b1;
27509: pixelout<=1'b0;
27510: pixelout<=1'b1;
27511: pixelout<=1'b1;
27512: pixelout<=1'b1;
27513: pixelout<=1'b1;
27514: pixelout<=1'b1;
27515: pixelout<=1'b1;
27516: pixelout<=1'b1;
27517: pixelout<=1'b1;
27518: pixelout<=1'b1;
27519: pixelout<=1'b0;
27520: pixelout<=1'b1;
27521: pixelout<=1'b0;
27522: pixelout<=1'b1;
27523: pixelout<=1'b1;
27524: pixelout<=1'b1;
27525: pixelout<=1'b0;
27526: pixelout<=1'b1;
27527: pixelout<=1'b1;
27528: pixelout<=1'b1;
27529: pixelout<=1'b1;
27530: pixelout<=1'b1;
27531: pixelout<=1'b1;
27532: pixelout<=1'b1;
27533: pixelout<=1'b1;
27534: pixelout<=1'b0;
27535: pixelout<=1'b1;
27536: pixelout<=1'b1;
27537: pixelout<=1'b1;
27538: pixelout<=1'b1;
27539: pixelout<=1'b1;
27540: pixelout<=1'b1;
27541: pixelout<=1'b1;
27542: pixelout<=1'b1;
27543: pixelout<=1'b1;
27544: pixelout<=1'b0;
27545: pixelout<=1'b1;
27546: pixelout<=1'b0;
27547: pixelout<=1'b1;
27548: pixelout<=1'b1;
27549: pixelout<=1'b1;
27550: pixelout<=1'b0;
27551: pixelout<=1'b1;
27552: pixelout<=1'b1;
27553: pixelout<=1'b1;
27554: pixelout<=1'b0;
27555: pixelout<=1'b1;
27556: pixelout<=1'b1;
27557: pixelout<=1'b1;
27558: pixelout<=1'b0;
27559: pixelout<=1'b1;
27560: pixelout<=1'b0;
27561: pixelout<=1'b1;
27562: pixelout<=1'b1;
27563: pixelout<=1'b1;
27564: pixelout<=1'b1;
27565: pixelout<=1'b1;
27566: pixelout<=1'b1;
27567: pixelout<=1'b1;
27568: pixelout<=1'b1;
27569: pixelout<=1'b1;
27570: pixelout<=1'b1;
27571: pixelout<=1'b0;
27572: pixelout<=1'b1;
27573: pixelout<=1'b0;
27574: pixelout<=1'b1;
27575: pixelout<=1'b1;
27576: pixelout<=1'b1;
27577: pixelout<=1'b0;
27578: pixelout<=1'b1;
27579: pixelout<=1'b1;
27580: pixelout<=1'b1;
27581: pixelout<=1'b1;
27582: pixelout<=1'b1;
27583: pixelout<=1'b1;
27584: pixelout<=1'b1;
27585: pixelout<=1'b1;
27586: pixelout<=1'b1;
27587: pixelout<=1'b1;
27588: pixelout<=1'b1;
27589: pixelout<=1'b1;
27590: pixelout<=1'b1;
27591: pixelout<=1'b1;
27592: pixelout<=1'b1;
27593: pixelout<=1'b1;
27594: pixelout<=1'b1;
27595: pixelout<=1'b1;
27596: pixelout<=1'b1;
27597: pixelout<=1'b1;
27598: pixelout<=1'b1;
27599: pixelout<=1'b1;
27600: pixelout<=1'b1;
27601: pixelout<=1'b1;
27602: pixelout<=1'b1;
27603: pixelout<=1'b1;
27604: pixelout<=1'b1;
27605: pixelout<=1'b1;
27606: pixelout<=1'b1;
27607: pixelout<=1'b1;
27608: pixelout<=1'b1;
27609: pixelout<=1'b1;
27610: pixelout<=1'b1;
27611: pixelout<=1'b1;
27612: pixelout<=1'b1;
27613: pixelout<=1'b1;
27614: pixelout<=1'b1;
27615: pixelout<=1'b1;
27616: pixelout<=1'b1;
27617: pixelout<=1'b1;
27618: pixelout<=1'b1;
27619: pixelout<=1'b0;
27620: pixelout<=1'b1;
27621: pixelout<=1'b1;
27622: pixelout<=1'b1;
27623: pixelout<=1'b1;
27624: pixelout<=1'b1;
27625: pixelout<=1'b0;
27626: pixelout<=1'b1;
27627: pixelout<=1'b1;
27628: pixelout<=1'b1;
27629: pixelout<=1'b1;
27630: pixelout<=1'b1;
27631: pixelout<=1'b1;
27632: pixelout<=1'b1;
27633: pixelout<=1'b1;
27634: pixelout<=1'b1;
27635: pixelout<=1'b0;
27636: pixelout<=1'b1;
27637: pixelout<=1'b0;
27638: pixelout<=1'b1;
27639: pixelout<=1'b1;
27640: pixelout<=1'b1;
27641: pixelout<=1'b0;
27642: pixelout<=1'b1;
27643: pixelout<=1'b0;
27644: pixelout<=1'b1;
27645: pixelout<=1'b1;
27646: pixelout<=1'b1;
27647: pixelout<=1'b1;
27648: pixelout<=1'b0;
27649: pixelout<=1'b1;
27650: pixelout<=1'b1;
27651: pixelout<=1'b1;
27652: pixelout<=1'b1;
27653: pixelout<=1'b1;
27654: pixelout<=1'b1;
27655: pixelout<=1'b1;
27656: pixelout<=1'b1;
27657: pixelout<=1'b1;
27658: pixelout<=1'b1;
27659: pixelout<=1'b1;
27660: pixelout<=1'b1;
27661: pixelout<=1'b0;
27662: pixelout<=1'b0;
27663: pixelout<=1'b1;
27664: pixelout<=1'b1;
27665: pixelout<=1'b1;
27666: pixelout<=1'b1;
27667: pixelout<=1'b0;
27668: pixelout<=1'b1;
27669: pixelout<=1'b1;
27670: pixelout<=1'b0;
27671: pixelout<=1'b1;
27672: pixelout<=1'b1;
27673: pixelout<=1'b1;
27674: pixelout<=1'b1;
27675: pixelout<=1'b1;
27676: pixelout<=1'b0;
27677: pixelout<=1'b1;
27678: pixelout<=1'b1;
27679: pixelout<=1'b1;
27680: pixelout<=1'b1;
27681: pixelout<=1'b1;
27682: pixelout<=1'b1;
27683: pixelout<=1'b1;
27684: pixelout<=1'b1;
27685: pixelout<=1'b1;
27686: pixelout<=1'b1;
27687: pixelout<=1'b0;
27688: pixelout<=1'b1;
27689: pixelout<=1'b0;
27690: pixelout<=1'b1;
27691: pixelout<=1'b1;
27692: pixelout<=1'b0;
27693: pixelout<=1'b1;
27694: pixelout<=1'b1;
27695: pixelout<=1'b1;
27696: pixelout<=1'b1;
27697: pixelout<=1'b1;
27698: pixelout<=1'b0;
27699: pixelout<=1'b1;
27700: pixelout<=1'b1;
27701: pixelout<=1'b1;
27702: pixelout<=1'b1;
27703: pixelout<=1'b1;
27704: pixelout<=1'b0;
27705: pixelout<=1'b0;
27706: pixelout<=1'b0;
27707: pixelout<=1'b0;
27708: pixelout<=1'b0;
27709: pixelout<=1'b1;
27710: pixelout<=1'b1;
27711: pixelout<=1'b1;
27712: pixelout<=1'b0;
27713: pixelout<=1'b1;
27714: pixelout<=1'b1;
27715: pixelout<=1'b1;
27716: pixelout<=1'b0;
27717: pixelout<=1'b1;
27718: pixelout<=1'b0;
27719: pixelout<=1'b1;
27720: pixelout<=1'b1;
27721: pixelout<=1'b1;
27722: pixelout<=1'b1;
27723: pixelout<=1'b0;
27724: pixelout<=1'b1;
27725: pixelout<=1'b1;
27726: pixelout<=1'b1;
27727: pixelout<=1'b1;
27728: pixelout<=1'b1;
27729: pixelout<=1'b1;
27730: pixelout<=1'b1;
27731: pixelout<=1'b1;
27732: pixelout<=1'b1;
27733: pixelout<=1'b1;
27734: pixelout<=1'b0;
27735: pixelout<=1'b1;
27736: pixelout<=1'b0;
27737: pixelout<=1'b1;
27738: pixelout<=1'b1;
27739: pixelout<=1'b0;
27740: pixelout<=1'b1;
27741: pixelout<=1'b1;
27742: pixelout<=1'b0;
27743: pixelout<=1'b1;
27744: pixelout<=1'b1;
27745: pixelout<=1'b1;
27746: pixelout<=1'b0;
27747: pixelout<=1'b1;
27748: pixelout<=1'b1;
27749: pixelout<=1'b0;
27750: pixelout<=1'b1;
27751: pixelout<=1'b1;
27752: pixelout<=1'b1;
27753: pixelout<=1'b1;
27754: pixelout<=1'b1;
27755: pixelout<=1'b1;
27756: pixelout<=1'b1;
27757: pixelout<=1'b1;
27758: pixelout<=1'b1;
27759: pixelout<=1'b0;
27760: pixelout<=1'b1;
27761: pixelout<=1'b0;
27762: pixelout<=1'b1;
27763: pixelout<=1'b1;
27764: pixelout<=1'b1;
27765: pixelout<=1'b0;
27766: pixelout<=1'b1;
27767: pixelout<=1'b1;
27768: pixelout<=1'b1;
27769: pixelout<=1'b1;
27770: pixelout<=1'b1;
27771: pixelout<=1'b1;
27772: pixelout<=1'b1;
27773: pixelout<=1'b1;
27774: pixelout<=1'b0;
27775: pixelout<=1'b1;
27776: pixelout<=1'b1;
27777: pixelout<=1'b1;
27778: pixelout<=1'b1;
27779: pixelout<=1'b1;
27780: pixelout<=1'b1;
27781: pixelout<=1'b1;
27782: pixelout<=1'b1;
27783: pixelout<=1'b1;
27784: pixelout<=1'b0;
27785: pixelout<=1'b1;
27786: pixelout<=1'b0;
27787: pixelout<=1'b1;
27788: pixelout<=1'b1;
27789: pixelout<=1'b1;
27790: pixelout<=1'b0;
27791: pixelout<=1'b1;
27792: pixelout<=1'b1;
27793: pixelout<=1'b1;
27794: pixelout<=1'b0;
27795: pixelout<=1'b1;
27796: pixelout<=1'b1;
27797: pixelout<=1'b1;
27798: pixelout<=1'b0;
27799: pixelout<=1'b1;
27800: pixelout<=1'b0;
27801: pixelout<=1'b1;
27802: pixelout<=1'b1;
27803: pixelout<=1'b1;
27804: pixelout<=1'b1;
27805: pixelout<=1'b1;
27806: pixelout<=1'b1;
27807: pixelout<=1'b1;
27808: pixelout<=1'b1;
27809: pixelout<=1'b1;
27810: pixelout<=1'b0;
27811: pixelout<=1'b1;
27812: pixelout<=1'b1;
27813: pixelout<=1'b0;
27814: pixelout<=1'b0;
27815: pixelout<=1'b0;
27816: pixelout<=1'b0;
27817: pixelout<=1'b0;
27818: pixelout<=1'b1;
27819: pixelout<=1'b1;
27820: pixelout<=1'b1;
27821: pixelout<=1'b1;
27822: pixelout<=1'b1;
27823: pixelout<=1'b1;
27824: pixelout<=1'b1;
27825: pixelout<=1'b1;
27826: pixelout<=1'b1;
27827: pixelout<=1'b1;
27828: pixelout<=1'b1;
27829: pixelout<=1'b1;
27830: pixelout<=1'b1;
27831: pixelout<=1'b1;
27832: pixelout<=1'b1;
27833: pixelout<=1'b1;
27834: pixelout<=1'b1;
27835: pixelout<=1'b1;
27836: pixelout<=1'b1;
27837: pixelout<=1'b1;
27838: pixelout<=1'b1;
27839: pixelout<=1'b1;
27840: pixelout<=1'b1;
27841: pixelout<=1'b1;
27842: pixelout<=1'b1;
27843: pixelout<=1'b1;
27844: pixelout<=1'b1;
27845: pixelout<=1'b1;
27846: pixelout<=1'b1;
27847: pixelout<=1'b1;
27848: pixelout<=1'b1;
27849: pixelout<=1'b1;
27850: pixelout<=1'b1;
27851: pixelout<=1'b1;
27852: pixelout<=1'b1;
27853: pixelout<=1'b1;
27854: pixelout<=1'b1;
27855: pixelout<=1'b1;
27856: pixelout<=1'b1;
27857: pixelout<=1'b1;
27858: pixelout<=1'b1;
27859: pixelout<=1'b0;
27860: pixelout<=1'b1;
27861: pixelout<=1'b1;
27862: pixelout<=1'b1;
27863: pixelout<=1'b0;
27864: pixelout<=1'b1;
27865: pixelout<=1'b0;
27866: pixelout<=1'b1;
27867: pixelout<=1'b1;
27868: pixelout<=1'b1;
27869: pixelout<=1'b1;
27870: pixelout<=1'b1;
27871: pixelout<=1'b1;
27872: pixelout<=1'b1;
27873: pixelout<=1'b1;
27874: pixelout<=1'b1;
27875: pixelout<=1'b0;
27876: pixelout<=1'b1;
27877: pixelout<=1'b0;
27878: pixelout<=1'b1;
27879: pixelout<=1'b1;
27880: pixelout<=1'b1;
27881: pixelout<=1'b0;
27882: pixelout<=1'b1;
27883: pixelout<=1'b0;
27884: pixelout<=1'b1;
27885: pixelout<=1'b1;
27886: pixelout<=1'b1;
27887: pixelout<=1'b1;
27888: pixelout<=1'b0;
27889: pixelout<=1'b1;
27890: pixelout<=1'b1;
27891: pixelout<=1'b0;
27892: pixelout<=1'b0;
27893: pixelout<=1'b1;
27894: pixelout<=1'b1;
27895: pixelout<=1'b1;
27896: pixelout<=1'b1;
27897: pixelout<=1'b1;
27898: pixelout<=1'b1;
27899: pixelout<=1'b1;
27900: pixelout<=1'b1;
27901: pixelout<=1'b1;
27902: pixelout<=1'b1;
27903: pixelout<=1'b0;
27904: pixelout<=1'b1;
27905: pixelout<=1'b1;
27906: pixelout<=1'b1;
27907: pixelout<=1'b0;
27908: pixelout<=1'b1;
27909: pixelout<=1'b1;
27910: pixelout<=1'b0;
27911: pixelout<=1'b1;
27912: pixelout<=1'b1;
27913: pixelout<=1'b1;
27914: pixelout<=1'b1;
27915: pixelout<=1'b1;
27916: pixelout<=1'b0;
27917: pixelout<=1'b1;
27918: pixelout<=1'b1;
27919: pixelout<=1'b1;
27920: pixelout<=1'b1;
27921: pixelout<=1'b1;
27922: pixelout<=1'b1;
27923: pixelout<=1'b1;
27924: pixelout<=1'b1;
27925: pixelout<=1'b1;
27926: pixelout<=1'b1;
27927: pixelout<=1'b0;
27928: pixelout<=1'b1;
27929: pixelout<=1'b0;
27930: pixelout<=1'b1;
27931: pixelout<=1'b1;
27932: pixelout<=1'b0;
27933: pixelout<=1'b1;
27934: pixelout<=1'b1;
27935: pixelout<=1'b1;
27936: pixelout<=1'b1;
27937: pixelout<=1'b1;
27938: pixelout<=1'b0;
27939: pixelout<=1'b1;
27940: pixelout<=1'b1;
27941: pixelout<=1'b1;
27942: pixelout<=1'b1;
27943: pixelout<=1'b1;
27944: pixelout<=1'b1;
27945: pixelout<=1'b1;
27946: pixelout<=1'b1;
27947: pixelout<=1'b1;
27948: pixelout<=1'b1;
27949: pixelout<=1'b1;
27950: pixelout<=1'b1;
27951: pixelout<=1'b1;
27952: pixelout<=1'b0;
27953: pixelout<=1'b1;
27954: pixelout<=1'b1;
27955: pixelout<=1'b1;
27956: pixelout<=1'b0;
27957: pixelout<=1'b1;
27958: pixelout<=1'b0;
27959: pixelout<=1'b1;
27960: pixelout<=1'b1;
27961: pixelout<=1'b1;
27962: pixelout<=1'b1;
27963: pixelout<=1'b0;
27964: pixelout<=1'b1;
27965: pixelout<=1'b1;
27966: pixelout<=1'b0;
27967: pixelout<=1'b0;
27968: pixelout<=1'b1;
27969: pixelout<=1'b1;
27970: pixelout<=1'b1;
27971: pixelout<=1'b1;
27972: pixelout<=1'b1;
27973: pixelout<=1'b1;
27974: pixelout<=1'b0;
27975: pixelout<=1'b1;
27976: pixelout<=1'b0;
27977: pixelout<=1'b1;
27978: pixelout<=1'b1;
27979: pixelout<=1'b0;
27980: pixelout<=1'b1;
27981: pixelout<=1'b1;
27982: pixelout<=1'b0;
27983: pixelout<=1'b1;
27984: pixelout<=1'b1;
27985: pixelout<=1'b0;
27986: pixelout<=1'b0;
27987: pixelout<=1'b1;
27988: pixelout<=1'b1;
27989: pixelout<=1'b0;
27990: pixelout<=1'b1;
27991: pixelout<=1'b1;
27992: pixelout<=1'b1;
27993: pixelout<=1'b1;
27994: pixelout<=1'b1;
27995: pixelout<=1'b1;
27996: pixelout<=1'b1;
27997: pixelout<=1'b1;
27998: pixelout<=1'b1;
27999: pixelout<=1'b0;
28000: pixelout<=1'b1;
28001: pixelout<=1'b0;
28002: pixelout<=1'b1;
28003: pixelout<=1'b1;
28004: pixelout<=1'b1;
28005: pixelout<=1'b0;
28006: pixelout<=1'b1;
28007: pixelout<=1'b0;
28008: pixelout<=1'b0;
28009: pixelout<=1'b1;
28010: pixelout<=1'b1;
28011: pixelout<=1'b1;
28012: pixelout<=1'b1;
28013: pixelout<=1'b1;
28014: pixelout<=1'b0;
28015: pixelout<=1'b1;
28016: pixelout<=1'b1;
28017: pixelout<=1'b0;
28018: pixelout<=1'b0;
28019: pixelout<=1'b1;
28020: pixelout<=1'b1;
28021: pixelout<=1'b1;
28022: pixelout<=1'b1;
28023: pixelout<=1'b1;
28024: pixelout<=1'b0;
28025: pixelout<=1'b1;
28026: pixelout<=1'b0;
28027: pixelout<=1'b1;
28028: pixelout<=1'b1;
28029: pixelout<=1'b1;
28030: pixelout<=1'b0;
28031: pixelout<=1'b1;
28032: pixelout<=1'b1;
28033: pixelout<=1'b1;
28034: pixelout<=1'b0;
28035: pixelout<=1'b1;
28036: pixelout<=1'b1;
28037: pixelout<=1'b1;
28038: pixelout<=1'b0;
28039: pixelout<=1'b1;
28040: pixelout<=1'b0;
28041: pixelout<=1'b1;
28042: pixelout<=1'b1;
28043: pixelout<=1'b0;
28044: pixelout<=1'b0;
28045: pixelout<=1'b1;
28046: pixelout<=1'b1;
28047: pixelout<=1'b1;
28048: pixelout<=1'b1;
28049: pixelout<=1'b1;
28050: pixelout<=1'b0;
28051: pixelout<=1'b1;
28052: pixelout<=1'b1;
28053: pixelout<=1'b0;
28054: pixelout<=1'b1;
28055: pixelout<=1'b1;
28056: pixelout<=1'b1;
28057: pixelout<=1'b1;
28058: pixelout<=1'b1;
28059: pixelout<=1'b1;
28060: pixelout<=1'b1;
28061: pixelout<=1'b1;
28062: pixelout<=1'b1;
28063: pixelout<=1'b1;
28064: pixelout<=1'b1;
28065: pixelout<=1'b1;
28066: pixelout<=1'b1;
28067: pixelout<=1'b1;
28068: pixelout<=1'b1;
28069: pixelout<=1'b1;
28070: pixelout<=1'b1;
28071: pixelout<=1'b1;
28072: pixelout<=1'b1;
28073: pixelout<=1'b1;
28074: pixelout<=1'b1;
28075: pixelout<=1'b1;
28076: pixelout<=1'b1;
28077: pixelout<=1'b1;
28078: pixelout<=1'b1;
28079: pixelout<=1'b1;
28080: pixelout<=1'b1;
28081: pixelout<=1'b1;
28082: pixelout<=1'b1;
28083: pixelout<=1'b1;
28084: pixelout<=1'b1;
28085: pixelout<=1'b1;
28086: pixelout<=1'b1;
28087: pixelout<=1'b1;
28088: pixelout<=1'b1;
28089: pixelout<=1'b1;
28090: pixelout<=1'b1;
28091: pixelout<=1'b1;
28092: pixelout<=1'b1;
28093: pixelout<=1'b1;
28094: pixelout<=1'b1;
28095: pixelout<=1'b1;
28096: pixelout<=1'b1;
28097: pixelout<=1'b1;
28098: pixelout<=1'b1;
28099: pixelout<=1'b1;
28100: pixelout<=1'b0;
28101: pixelout<=1'b0;
28102: pixelout<=1'b0;
28103: pixelout<=1'b1;
28104: pixelout<=1'b1;
28105: pixelout<=1'b1;
28106: pixelout<=1'b0;
28107: pixelout<=1'b0;
28108: pixelout<=1'b0;
28109: pixelout<=1'b1;
28110: pixelout<=1'b1;
28111: pixelout<=1'b1;
28112: pixelout<=1'b1;
28113: pixelout<=1'b1;
28114: pixelout<=1'b1;
28115: pixelout<=1'b0;
28116: pixelout<=1'b1;
28117: pixelout<=1'b1;
28118: pixelout<=1'b0;
28119: pixelout<=1'b0;
28120: pixelout<=1'b0;
28121: pixelout<=1'b0;
28122: pixelout<=1'b1;
28123: pixelout<=1'b0;
28124: pixelout<=1'b1;
28125: pixelout<=1'b1;
28126: pixelout<=1'b1;
28127: pixelout<=1'b1;
28128: pixelout<=1'b1;
28129: pixelout<=1'b0;
28130: pixelout<=1'b0;
28131: pixelout<=1'b1;
28132: pixelout<=1'b1;
28133: pixelout<=1'b1;
28134: pixelout<=1'b1;
28135: pixelout<=1'b1;
28136: pixelout<=1'b0;
28137: pixelout<=1'b0;
28138: pixelout<=1'b0;
28139: pixelout<=1'b1;
28140: pixelout<=1'b0;
28141: pixelout<=1'b0;
28142: pixelout<=1'b0;
28143: pixelout<=1'b0;
28144: pixelout<=1'b1;
28145: pixelout<=1'b1;
28146: pixelout<=1'b1;
28147: pixelout<=1'b0;
28148: pixelout<=1'b1;
28149: pixelout<=1'b1;
28150: pixelout<=1'b0;
28151: pixelout<=1'b1;
28152: pixelout<=1'b1;
28153: pixelout<=1'b1;
28154: pixelout<=1'b1;
28155: pixelout<=1'b1;
28156: pixelout<=1'b1;
28157: pixelout<=1'b0;
28158: pixelout<=1'b0;
28159: pixelout<=1'b0;
28160: pixelout<=1'b0;
28161: pixelout<=1'b1;
28162: pixelout<=1'b1;
28163: pixelout<=1'b1;
28164: pixelout<=1'b0;
28165: pixelout<=1'b0;
28166: pixelout<=1'b0;
28167: pixelout<=1'b1;
28168: pixelout<=1'b1;
28169: pixelout<=1'b1;
28170: pixelout<=1'b0;
28171: pixelout<=1'b0;
28172: pixelout<=1'b1;
28173: pixelout<=1'b0;
28174: pixelout<=1'b1;
28175: pixelout<=1'b1;
28176: pixelout<=1'b1;
28177: pixelout<=1'b1;
28178: pixelout<=1'b0;
28179: pixelout<=1'b1;
28180: pixelout<=1'b1;
28181: pixelout<=1'b1;
28182: pixelout<=1'b1;
28183: pixelout<=1'b1;
28184: pixelout<=1'b1;
28185: pixelout<=1'b0;
28186: pixelout<=1'b0;
28187: pixelout<=1'b0;
28188: pixelout<=1'b0;
28189: pixelout<=1'b1;
28190: pixelout<=1'b1;
28191: pixelout<=1'b1;
28192: pixelout<=1'b1;
28193: pixelout<=1'b0;
28194: pixelout<=1'b0;
28195: pixelout<=1'b0;
28196: pixelout<=1'b0;
28197: pixelout<=1'b1;
28198: pixelout<=1'b0;
28199: pixelout<=1'b1;
28200: pixelout<=1'b1;
28201: pixelout<=1'b1;
28202: pixelout<=1'b1;
28203: pixelout<=1'b1;
28204: pixelout<=1'b0;
28205: pixelout<=1'b0;
28206: pixelout<=1'b1;
28207: pixelout<=1'b1;
28208: pixelout<=1'b1;
28209: pixelout<=1'b1;
28210: pixelout<=1'b1;
28211: pixelout<=1'b0;
28212: pixelout<=1'b0;
28213: pixelout<=1'b0;
28214: pixelout<=1'b0;
28215: pixelout<=1'b1;
28216: pixelout<=1'b1;
28217: pixelout<=1'b0;
28218: pixelout<=1'b0;
28219: pixelout<=1'b1;
28220: pixelout<=1'b0;
28221: pixelout<=1'b1;
28222: pixelout<=1'b1;
28223: pixelout<=1'b0;
28224: pixelout<=1'b0;
28225: pixelout<=1'b1;
28226: pixelout<=1'b0;
28227: pixelout<=1'b1;
28228: pixelout<=1'b1;
28229: pixelout<=1'b0;
28230: pixelout<=1'b0;
28231: pixelout<=1'b0;
28232: pixelout<=1'b1;
28233: pixelout<=1'b1;
28234: pixelout<=1'b1;
28235: pixelout<=1'b1;
28236: pixelout<=1'b1;
28237: pixelout<=1'b1;
28238: pixelout<=1'b1;
28239: pixelout<=1'b0;
28240: pixelout<=1'b1;
28241: pixelout<=1'b1;
28242: pixelout<=1'b0;
28243: pixelout<=1'b0;
28244: pixelout<=1'b0;
28245: pixelout<=1'b0;
28246: pixelout<=1'b1;
28247: pixelout<=1'b0;
28248: pixelout<=1'b0;
28249: pixelout<=1'b1;
28250: pixelout<=1'b1;
28251: pixelout<=1'b1;
28252: pixelout<=1'b1;
28253: pixelout<=1'b1;
28254: pixelout<=1'b1;
28255: pixelout<=1'b0;
28256: pixelout<=1'b0;
28257: pixelout<=1'b1;
28258: pixelout<=1'b1;
28259: pixelout<=1'b1;
28260: pixelout<=1'b1;
28261: pixelout<=1'b1;
28262: pixelout<=1'b1;
28263: pixelout<=1'b1;
28264: pixelout<=1'b0;
28265: pixelout<=1'b1;
28266: pixelout<=1'b1;
28267: pixelout<=1'b0;
28268: pixelout<=1'b0;
28269: pixelout<=1'b0;
28270: pixelout<=1'b0;
28271: pixelout<=1'b1;
28272: pixelout<=1'b1;
28273: pixelout<=1'b1;
28274: pixelout<=1'b0;
28275: pixelout<=1'b1;
28276: pixelout<=1'b1;
28277: pixelout<=1'b1;
28278: pixelout<=1'b0;
28279: pixelout<=1'b1;
28280: pixelout<=1'b1;
28281: pixelout<=1'b0;
28282: pixelout<=1'b0;
28283: pixelout<=1'b1;
28284: pixelout<=1'b1;
28285: pixelout<=1'b1;
28286: pixelout<=1'b1;
28287: pixelout<=1'b1;
28288: pixelout<=1'b1;
28289: pixelout<=1'b0;
28290: pixelout<=1'b1;
28291: pixelout<=1'b1;
28292: pixelout<=1'b1;
28293: pixelout<=1'b1;
28294: pixelout<=1'b0;
28295: pixelout<=1'b0;
28296: pixelout<=1'b0;
28297: pixelout<=1'b0;
28298: pixelout<=1'b1;
28299: pixelout<=1'b1;
28300: pixelout<=1'b1;
28301: pixelout<=1'b1;
28302: pixelout<=1'b1;
28303: pixelout<=1'b1;
28304: pixelout<=1'b1;
28305: pixelout<=1'b1;
28306: pixelout<=1'b1;
28307: pixelout<=1'b1;
28308: pixelout<=1'b1;
28309: pixelout<=1'b1;
28310: pixelout<=1'b1;
28311: pixelout<=1'b1;
28312: pixelout<=1'b1;
28313: pixelout<=1'b1;
28314: pixelout<=1'b1;
28315: pixelout<=1'b1;
28316: pixelout<=1'b1;
28317: pixelout<=1'b1;
28318: pixelout<=1'b1;
28319: pixelout<=1'b1;
28320: pixelout<=1'b1;
28321: pixelout<=1'b1;
28322: pixelout<=1'b1;
28323: pixelout<=1'b1;
28324: pixelout<=1'b1;
28325: pixelout<=1'b1;
28326: pixelout<=1'b1;
28327: pixelout<=1'b1;
28328: pixelout<=1'b1;
28329: pixelout<=1'b1;
28330: pixelout<=1'b1;
28331: pixelout<=1'b1;
28332: pixelout<=1'b1;
28333: pixelout<=1'b1;
28334: pixelout<=1'b1;
28335: pixelout<=1'b1;
28336: pixelout<=1'b1;
28337: pixelout<=1'b1;
28338: pixelout<=1'b1;
28339: pixelout<=1'b1;
28340: pixelout<=1'b1;
28341: pixelout<=1'b1;
28342: pixelout<=1'b1;
28343: pixelout<=1'b1;
28344: pixelout<=1'b1;
28345: pixelout<=1'b1;
28346: pixelout<=1'b1;
28347: pixelout<=1'b1;
28348: pixelout<=1'b1;
28349: pixelout<=1'b1;
28350: pixelout<=1'b1;
28351: pixelout<=1'b1;
28352: pixelout<=1'b1;
28353: pixelout<=1'b1;
28354: pixelout<=1'b1;
28355: pixelout<=1'b1;
28356: pixelout<=1'b1;
28357: pixelout<=1'b1;
28358: pixelout<=1'b1;
28359: pixelout<=1'b1;
28360: pixelout<=1'b1;
28361: pixelout<=1'b0;
28362: pixelout<=1'b1;
28363: pixelout<=1'b1;
28364: pixelout<=1'b1;
28365: pixelout<=1'b1;
28366: pixelout<=1'b1;
28367: pixelout<=1'b1;
28368: pixelout<=1'b1;
28369: pixelout<=1'b1;
28370: pixelout<=1'b1;
28371: pixelout<=1'b1;
28372: pixelout<=1'b1;
28373: pixelout<=1'b1;
28374: pixelout<=1'b1;
28375: pixelout<=1'b1;
28376: pixelout<=1'b1;
28377: pixelout<=1'b1;
28378: pixelout<=1'b1;
28379: pixelout<=1'b1;
28380: pixelout<=1'b1;
28381: pixelout<=1'b1;
28382: pixelout<=1'b1;
28383: pixelout<=1'b1;
28384: pixelout<=1'b1;
28385: pixelout<=1'b1;
28386: pixelout<=1'b1;
28387: pixelout<=1'b1;
28388: pixelout<=1'b1;
28389: pixelout<=1'b1;
28390: pixelout<=1'b1;
28391: pixelout<=1'b1;
28392: pixelout<=1'b1;
28393: pixelout<=1'b1;
28394: pixelout<=1'b1;
28395: pixelout<=1'b1;
28396: pixelout<=1'b1;
28397: pixelout<=1'b1;
28398: pixelout<=1'b1;
28399: pixelout<=1'b1;
28400: pixelout<=1'b1;
28401: pixelout<=1'b1;
28402: pixelout<=1'b1;
28403: pixelout<=1'b1;
28404: pixelout<=1'b1;
28405: pixelout<=1'b1;
28406: pixelout<=1'b1;
28407: pixelout<=1'b1;
28408: pixelout<=1'b1;
28409: pixelout<=1'b1;
28410: pixelout<=1'b1;
28411: pixelout<=1'b1;
28412: pixelout<=1'b1;
28413: pixelout<=1'b1;
28414: pixelout<=1'b1;
28415: pixelout<=1'b1;
28416: pixelout<=1'b1;
28417: pixelout<=1'b1;
28418: pixelout<=1'b1;
28419: pixelout<=1'b1;
28420: pixelout<=1'b1;
28421: pixelout<=1'b1;
28422: pixelout<=1'b1;
28423: pixelout<=1'b1;
28424: pixelout<=1'b1;
28425: pixelout<=1'b1;
28426: pixelout<=1'b1;
28427: pixelout<=1'b1;
28428: pixelout<=1'b1;
28429: pixelout<=1'b1;
28430: pixelout<=1'b1;
28431: pixelout<=1'b1;
28432: pixelout<=1'b1;
28433: pixelout<=1'b1;
28434: pixelout<=1'b1;
28435: pixelout<=1'b1;
28436: pixelout<=1'b0;
28437: pixelout<=1'b1;
28438: pixelout<=1'b1;
28439: pixelout<=1'b1;
28440: pixelout<=1'b1;
28441: pixelout<=1'b1;
28442: pixelout<=1'b1;
28443: pixelout<=1'b1;
28444: pixelout<=1'b1;
28445: pixelout<=1'b1;
28446: pixelout<=1'b1;
28447: pixelout<=1'b1;
28448: pixelout<=1'b1;
28449: pixelout<=1'b1;
28450: pixelout<=1'b1;
28451: pixelout<=1'b1;
28452: pixelout<=1'b1;
28453: pixelout<=1'b1;
28454: pixelout<=1'b1;
28455: pixelout<=1'b1;
28456: pixelout<=1'b1;
28457: pixelout<=1'b1;
28458: pixelout<=1'b1;
28459: pixelout<=1'b1;
28460: pixelout<=1'b1;
28461: pixelout<=1'b1;
28462: pixelout<=1'b1;
28463: pixelout<=1'b1;
28464: pixelout<=1'b1;
28465: pixelout<=1'b1;
28466: pixelout<=1'b1;
28467: pixelout<=1'b1;
28468: pixelout<=1'b1;
28469: pixelout<=1'b1;
28470: pixelout<=1'b1;
28471: pixelout<=1'b1;
28472: pixelout<=1'b1;
28473: pixelout<=1'b1;
28474: pixelout<=1'b1;
28475: pixelout<=1'b1;
28476: pixelout<=1'b1;
28477: pixelout<=1'b1;
28478: pixelout<=1'b1;
28479: pixelout<=1'b1;
28480: pixelout<=1'b1;
28481: pixelout<=1'b1;
28482: pixelout<=1'b1;
28483: pixelout<=1'b1;
28484: pixelout<=1'b1;
28485: pixelout<=1'b0;
28486: pixelout<=1'b1;
28487: pixelout<=1'b1;
28488: pixelout<=1'b0;
28489: pixelout<=1'b1;
28490: pixelout<=1'b1;
28491: pixelout<=1'b1;
28492: pixelout<=1'b1;
28493: pixelout<=1'b1;
28494: pixelout<=1'b1;
28495: pixelout<=1'b1;
28496: pixelout<=1'b1;
28497: pixelout<=1'b1;
28498: pixelout<=1'b1;
28499: pixelout<=1'b1;
28500: pixelout<=1'b1;
28501: pixelout<=1'b1;
28502: pixelout<=1'b1;
28503: pixelout<=1'b1;
28504: pixelout<=1'b1;
28505: pixelout<=1'b1;
28506: pixelout<=1'b1;
28507: pixelout<=1'b1;
28508: pixelout<=1'b1;
28509: pixelout<=1'b1;
28510: pixelout<=1'b1;
28511: pixelout<=1'b1;
28512: pixelout<=1'b1;
28513: pixelout<=1'b1;
28514: pixelout<=1'b1;
28515: pixelout<=1'b1;
28516: pixelout<=1'b1;
28517: pixelout<=1'b1;
28518: pixelout<=1'b1;
28519: pixelout<=1'b1;
28520: pixelout<=1'b1;
28521: pixelout<=1'b1;
28522: pixelout<=1'b1;
28523: pixelout<=1'b1;
28524: pixelout<=1'b1;
28525: pixelout<=1'b1;
28526: pixelout<=1'b1;
28527: pixelout<=1'b1;
28528: pixelout<=1'b1;
28529: pixelout<=1'b1;
28530: pixelout<=1'b1;
28531: pixelout<=1'b1;
28532: pixelout<=1'b1;
28533: pixelout<=1'b1;
28534: pixelout<=1'b1;
28535: pixelout<=1'b1;
28536: pixelout<=1'b1;
28537: pixelout<=1'b1;
28538: pixelout<=1'b1;
28539: pixelout<=1'b1;
28540: pixelout<=1'b1;
28541: pixelout<=1'b1;
28542: pixelout<=1'b1;
28543: pixelout<=1'b1;
28544: pixelout<=1'b1;
28545: pixelout<=1'b1;
28546: pixelout<=1'b1;
28547: pixelout<=1'b1;
28548: pixelout<=1'b1;
28549: pixelout<=1'b1;
28550: pixelout<=1'b1;
28551: pixelout<=1'b1;
28552: pixelout<=1'b1;
28553: pixelout<=1'b1;
28554: pixelout<=1'b1;
28555: pixelout<=1'b1;
28556: pixelout<=1'b1;
28557: pixelout<=1'b1;
28558: pixelout<=1'b1;
28559: pixelout<=1'b1;
28560: pixelout<=1'b1;
28561: pixelout<=1'b1;
28562: pixelout<=1'b1;
28563: pixelout<=1'b1;
28564: pixelout<=1'b1;
28565: pixelout<=1'b1;
28566: pixelout<=1'b1;
28567: pixelout<=1'b1;
28568: pixelout<=1'b1;
28569: pixelout<=1'b1;
28570: pixelout<=1'b1;
28571: pixelout<=1'b1;
28572: pixelout<=1'b1;
28573: pixelout<=1'b1;
28574: pixelout<=1'b1;
28575: pixelout<=1'b1;
28576: pixelout<=1'b1;
28577: pixelout<=1'b1;
28578: pixelout<=1'b1;
28579: pixelout<=1'b1;
28580: pixelout<=1'b1;
28581: pixelout<=1'b1;
28582: pixelout<=1'b1;
28583: pixelout<=1'b1;
28584: pixelout<=1'b1;
28585: pixelout<=1'b1;
28586: pixelout<=1'b1;
28587: pixelout<=1'b1;
28588: pixelout<=1'b1;
28589: pixelout<=1'b1;
28590: pixelout<=1'b1;
28591: pixelout<=1'b1;
28592: pixelout<=1'b1;
28593: pixelout<=1'b1;
28594: pixelout<=1'b1;
28595: pixelout<=1'b1;
28596: pixelout<=1'b1;
28597: pixelout<=1'b1;
28598: pixelout<=1'b0;
28599: pixelout<=1'b0;
28600: pixelout<=1'b0;
28601: pixelout<=1'b1;
28602: pixelout<=1'b1;
28603: pixelout<=1'b1;
28604: pixelout<=1'b1;
28605: pixelout<=1'b1;
28606: pixelout<=1'b1;
28607: pixelout<=1'b1;
28608: pixelout<=1'b1;
28609: pixelout<=1'b1;
28610: pixelout<=1'b1;
28611: pixelout<=1'b1;
28612: pixelout<=1'b1;
28613: pixelout<=1'b1;
28614: pixelout<=1'b1;
28615: pixelout<=1'b1;
28616: pixelout<=1'b1;
28617: pixelout<=1'b1;
28618: pixelout<=1'b1;
28619: pixelout<=1'b1;
28620: pixelout<=1'b1;
28621: pixelout<=1'b1;
28622: pixelout<=1'b1;
28623: pixelout<=1'b1;
28624: pixelout<=1'b1;
28625: pixelout<=1'b1;
28626: pixelout<=1'b1;
28627: pixelout<=1'b1;
28628: pixelout<=1'b1;
28629: pixelout<=1'b1;
28630: pixelout<=1'b1;
28631: pixelout<=1'b1;
28632: pixelout<=1'b1;
28633: pixelout<=1'b1;
28634: pixelout<=1'b1;
28635: pixelout<=1'b1;
28636: pixelout<=1'b0;
28637: pixelout<=1'b0;
28638: pixelout<=1'b0;
28639: pixelout<=1'b0;
28640: pixelout<=1'b1;
28641: pixelout<=1'b1;
28642: pixelout<=1'b1;
28643: pixelout<=1'b1;
28644: pixelout<=1'b1;
28645: pixelout<=1'b1;
28646: pixelout<=1'b1;
28647: pixelout<=1'b1;
28648: pixelout<=1'b1;
28649: pixelout<=1'b1;
28650: pixelout<=1'b1;
28651: pixelout<=1'b1;
28652: pixelout<=1'b1;
28653: pixelout<=1'b1;
28654: pixelout<=1'b1;
28655: pixelout<=1'b1;
28656: pixelout<=1'b1;
28657: pixelout<=1'b1;
28658: pixelout<=1'b1;
28659: pixelout<=1'b1;
28660: pixelout<=1'b1;
28661: pixelout<=1'b1;
28662: pixelout<=1'b1;
28663: pixelout<=1'b1;
28664: pixelout<=1'b1;
28665: pixelout<=1'b1;
28666: pixelout<=1'b1;
28667: pixelout<=1'b1;
28668: pixelout<=1'b1;
28669: pixelout<=1'b1;
28670: pixelout<=1'b1;
28671: pixelout<=1'b1;
28672: pixelout<=1'b1;
28673: pixelout<=1'b0;
28674: pixelout<=1'b0;
28675: pixelout<=1'b0;
28676: pixelout<=1'b1;
28677: pixelout<=1'b1;
28678: pixelout<=1'b1;
28679: pixelout<=1'b1;
28680: pixelout<=1'b1;
28681: pixelout<=1'b1;
28682: pixelout<=1'b1;
28683: pixelout<=1'b1;
28684: pixelout<=1'b1;
28685: pixelout<=1'b1;
28686: pixelout<=1'b1;
28687: pixelout<=1'b1;
28688: pixelout<=1'b1;
28689: pixelout<=1'b1;
28690: pixelout<=1'b1;
28691: pixelout<=1'b1;
28692: pixelout<=1'b1;
28693: pixelout<=1'b1;
28694: pixelout<=1'b1;
28695: pixelout<=1'b1;
28696: pixelout<=1'b1;
28697: pixelout<=1'b1;
28698: pixelout<=1'b1;
28699: pixelout<=1'b1;
28700: pixelout<=1'b1;
28701: pixelout<=1'b1;
28702: pixelout<=1'b1;
28703: pixelout<=1'b1;
28704: pixelout<=1'b1;
28705: pixelout<=1'b1;
28706: pixelout<=1'b1;
28707: pixelout<=1'b1;
28708: pixelout<=1'b1;
28709: pixelout<=1'b1;
28710: pixelout<=1'b1;
28711: pixelout<=1'b1;
28712: pixelout<=1'b1;
28713: pixelout<=1'b1;
28714: pixelout<=1'b1;
28715: pixelout<=1'b1;
28716: pixelout<=1'b1;
28717: pixelout<=1'b1;
28718: pixelout<=1'b1;
28719: pixelout<=1'b1;
28720: pixelout<=1'b1;
28721: pixelout<=1'b1;
28722: pixelout<=1'b0;
28723: pixelout<=1'b0;
28724: pixelout<=1'b0;
28725: pixelout<=1'b1;
28726: pixelout<=1'b1;
28727: pixelout<=1'b0;
28728: pixelout<=1'b1;
28729: pixelout<=1'b1;
28730: pixelout<=1'b1;
28731: pixelout<=1'b1;
28732: pixelout<=1'b1;
28733: pixelout<=1'b1;
28734: pixelout<=1'b1;
28735: pixelout<=1'b1;
28736: pixelout<=1'b1;
28737: pixelout<=1'b1;
28738: pixelout<=1'b1;
28739: pixelout<=1'b1;
28740: pixelout<=1'b1;
28741: pixelout<=1'b1;
28742: pixelout<=1'b1;
28743: pixelout<=1'b1;
28744: pixelout<=1'b1;
28745: pixelout<=1'b1;
28746: pixelout<=1'b1;
28747: pixelout<=1'b1;
28748: pixelout<=1'b1;
28749: pixelout<=1'b1;
28750: pixelout<=1'b1;
28751: pixelout<=1'b1;
28752: pixelout<=1'b1;
28753: pixelout<=1'b1;
28754: pixelout<=1'b1;
28755: pixelout<=1'b1;
28756: pixelout<=1'b1;
28757: pixelout<=1'b1;
28758: pixelout<=1'b1;
28759: pixelout<=1'b1;
28760: pixelout<=1'b1;
28761: pixelout<=1'b1;
28762: pixelout<=1'b1;
28763: pixelout<=1'b1;
28764: pixelout<=1'b1;
28765: pixelout<=1'b1;
28766: pixelout<=1'b1;
28767: pixelout<=1'b1;
28768: pixelout<=1'b1;
28769: pixelout<=1'b1;
28770: pixelout<=1'b1;
28771: pixelout<=1'b1;
28772: pixelout<=1'b1;
28773: pixelout<=1'b1;
28774: pixelout<=1'b1;
28775: pixelout<=1'b1;
28776: pixelout<=1'b1;
28777: pixelout<=1'b1;
28778: pixelout<=1'b1;
28779: pixelout<=1'b1;
28780: pixelout<=1'b1;
28781: pixelout<=1'b1;
28782: pixelout<=1'b1;
28783: pixelout<=1'b1;
28784: pixelout<=1'b1;
28785: pixelout<=1'b1;
28786: pixelout<=1'b1;
28787: pixelout<=1'b1;
28788: pixelout<=1'b1;
28789: pixelout<=1'b1;
28790: pixelout<=1'b1;
28791: pixelout<=1'b1;
28792: pixelout<=1'b1;
28793: pixelout<=1'b1;
28794: pixelout<=1'b1;
28795: pixelout<=1'b1;
28796: pixelout<=1'b1;
28797: pixelout<=1'b1;
28798: pixelout<=1'b1;
28799: pixelout<=1'b1;
28800: pixelout<=1'b1;
28801: pixelout<=1'b1;
28802: pixelout<=1'b1;
28803: pixelout<=1'b1;
28804: pixelout<=1'b1;
28805: pixelout<=1'b1;
28806: pixelout<=1'b1;
28807: pixelout<=1'b1;
28808: pixelout<=1'b1;
28809: pixelout<=1'b1;
28810: pixelout<=1'b1;
28811: pixelout<=1'b1;
28812: pixelout<=1'b1;
28813: pixelout<=1'b1;
28814: pixelout<=1'b1;
28815: pixelout<=1'b1;
28816: pixelout<=1'b1;
28817: pixelout<=1'b1;
28818: pixelout<=1'b1;
28819: pixelout<=1'b1;
28820: pixelout<=1'b1;
28821: pixelout<=1'b1;
28822: pixelout<=1'b1;
28823: pixelout<=1'b1;
28824: pixelout<=1'b1;
28825: pixelout<=1'b1;
28826: pixelout<=1'b1;
28827: pixelout<=1'b1;
28828: pixelout<=1'b1;
28829: pixelout<=1'b1;
28830: pixelout<=1'b1;
28831: pixelout<=1'b1;
28832: pixelout<=1'b1;
28833: pixelout<=1'b1;
28834: pixelout<=1'b1;
28835: pixelout<=1'b1;
28836: pixelout<=1'b1;
28837: pixelout<=1'b1;
28838: pixelout<=1'b1;
28839: pixelout<=1'b1;
28840: pixelout<=1'b1;
28841: pixelout<=1'b1;
28842: pixelout<=1'b1;
28843: pixelout<=1'b1;
28844: pixelout<=1'b1;
28845: pixelout<=1'b1;
28846: pixelout<=1'b1;
28847: pixelout<=1'b1;
28848: pixelout<=1'b1;
28849: pixelout<=1'b1;
28850: pixelout<=1'b1;
28851: pixelout<=1'b1;
28852: pixelout<=1'b1;
28853: pixelout<=1'b1;
28854: pixelout<=1'b1;
28855: pixelout<=1'b1;
28856: pixelout<=1'b1;
28857: pixelout<=1'b1;
28858: pixelout<=1'b1;
28859: pixelout<=1'b1;
28860: pixelout<=1'b1;
28861: pixelout<=1'b1;
28862: pixelout<=1'b1;
28863: pixelout<=1'b1;
28864: pixelout<=1'b1;
28865: pixelout<=1'b1;
28866: pixelout<=1'b1;
28867: pixelout<=1'b1;
28868: pixelout<=1'b1;
28869: pixelout<=1'b1;
28870: pixelout<=1'b1;
28871: pixelout<=1'b1;
28872: pixelout<=1'b1;
28873: pixelout<=1'b1;
28874: pixelout<=1'b1;
28875: pixelout<=1'b1;
28876: pixelout<=1'b1;
28877: pixelout<=1'b1;
28878: pixelout<=1'b1;
28879: pixelout<=1'b1;
28880: pixelout<=1'b1;
28881: pixelout<=1'b1;
28882: pixelout<=1'b1;
28883: pixelout<=1'b1;
28884: pixelout<=1'b1;
28885: pixelout<=1'b1;
28886: pixelout<=1'b1;
28887: pixelout<=1'b1;
28888: pixelout<=1'b1;
28889: pixelout<=1'b1;
28890: pixelout<=1'b1;
28891: pixelout<=1'b1;
28892: pixelout<=1'b1;
28893: pixelout<=1'b1;
28894: pixelout<=1'b1;
28895: pixelout<=1'b1;
28896: pixelout<=1'b1;
28897: pixelout<=1'b1;
28898: pixelout<=1'b1;
28899: pixelout<=1'b1;
28900: pixelout<=1'b1;
28901: pixelout<=1'b1;
28902: pixelout<=1'b1;
28903: pixelout<=1'b1;
28904: pixelout<=1'b1;
28905: pixelout<=1'b1;
28906: pixelout<=1'b1;
28907: pixelout<=1'b1;
28908: pixelout<=1'b1;
28909: pixelout<=1'b1;
28910: pixelout<=1'b1;
28911: pixelout<=1'b1;
28912: pixelout<=1'b1;
28913: pixelout<=1'b1;
28914: pixelout<=1'b1;
28915: pixelout<=1'b1;
28916: pixelout<=1'b1;
28917: pixelout<=1'b1;
28918: pixelout<=1'b1;
28919: pixelout<=1'b1;
28920: pixelout<=1'b1;
28921: pixelout<=1'b1;
28922: pixelout<=1'b1;
28923: pixelout<=1'b1;
28924: pixelout<=1'b1;
28925: pixelout<=1'b1;
28926: pixelout<=1'b1;
28927: pixelout<=1'b1;
28928: pixelout<=1'b1;
28929: pixelout<=1'b1;
28930: pixelout<=1'b1;
28931: pixelout<=1'b1;
28932: pixelout<=1'b1;
28933: pixelout<=1'b1;
28934: pixelout<=1'b1;
28935: pixelout<=1'b1;
28936: pixelout<=1'b1;
28937: pixelout<=1'b1;
28938: pixelout<=1'b1;
28939: pixelout<=1'b1;
28940: pixelout<=1'b1;
28941: pixelout<=1'b1;
28942: pixelout<=1'b1;
28943: pixelout<=1'b1;
28944: pixelout<=1'b1;
28945: pixelout<=1'b1;
28946: pixelout<=1'b1;
28947: pixelout<=1'b1;
28948: pixelout<=1'b1;
28949: pixelout<=1'b1;
28950: pixelout<=1'b1;
28951: pixelout<=1'b1;
28952: pixelout<=1'b1;
28953: pixelout<=1'b1;
28954: pixelout<=1'b1;
28955: pixelout<=1'b1;
28956: pixelout<=1'b1;
28957: pixelout<=1'b1;
28958: pixelout<=1'b1;
28959: pixelout<=1'b1;
28960: pixelout<=1'b1;
28961: pixelout<=1'b1;
28962: pixelout<=1'b1;
28963: pixelout<=1'b1;
28964: pixelout<=1'b1;
28965: pixelout<=1'b1;
28966: pixelout<=1'b1;
28967: pixelout<=1'b1;
28968: pixelout<=1'b1;
28969: pixelout<=1'b1;
28970: pixelout<=1'b1;
28971: pixelout<=1'b1;
28972: pixelout<=1'b1;
28973: pixelout<=1'b1;
28974: pixelout<=1'b1;
28975: pixelout<=1'b1;
28976: pixelout<=1'b1;
28977: pixelout<=1'b1;
28978: pixelout<=1'b1;
28979: pixelout<=1'b1;
28980: pixelout<=1'b1;
28981: pixelout<=1'b1;
28982: pixelout<=1'b1;
28983: pixelout<=1'b1;
28984: pixelout<=1'b1;
28985: pixelout<=1'b1;
28986: pixelout<=1'b1;
28987: pixelout<=1'b1;
28988: pixelout<=1'b1;
28989: pixelout<=1'b1;
28990: pixelout<=1'b1;
28991: pixelout<=1'b1;
28992: pixelout<=1'b1;
28993: pixelout<=1'b1;
28994: pixelout<=1'b1;
28995: pixelout<=1'b1;
28996: pixelout<=1'b1;
28997: pixelout<=1'b1;
28998: pixelout<=1'b1;
28999: pixelout<=1'b1;
29000: pixelout<=1'b1;
29001: pixelout<=1'b1;
29002: pixelout<=1'b1;
29003: pixelout<=1'b1;
29004: pixelout<=1'b1;
29005: pixelout<=1'b1;
29006: pixelout<=1'b1;
29007: pixelout<=1'b1;
29008: pixelout<=1'b1;
29009: pixelout<=1'b1;
29010: pixelout<=1'b1;
29011: pixelout<=1'b1;
29012: pixelout<=1'b1;
29013: pixelout<=1'b1;
29014: pixelout<=1'b1;
29015: pixelout<=1'b1;
29016: pixelout<=1'b1;
29017: pixelout<=1'b1;
29018: pixelout<=1'b1;
29019: pixelout<=1'b1;
29020: pixelout<=1'b1;
29021: pixelout<=1'b1;
29022: pixelout<=1'b1;
29023: pixelout<=1'b1;
29024: pixelout<=1'b1;
29025: pixelout<=1'b1;
29026: pixelout<=1'b1;
29027: pixelout<=1'b1;
29028: pixelout<=1'b1;
29029: pixelout<=1'b1;
29030: pixelout<=1'b1;
29031: pixelout<=1'b1;
29032: pixelout<=1'b1;
29033: pixelout<=1'b1;
29034: pixelout<=1'b1;
29035: pixelout<=1'b1;
29036: pixelout<=1'b1;
29037: pixelout<=1'b1;
29038: pixelout<=1'b1;
29039: pixelout<=1'b1;
29040: pixelout<=1'b1;
29041: pixelout<=1'b1;
29042: pixelout<=1'b1;
29043: pixelout<=1'b1;
29044: pixelout<=1'b1;
29045: pixelout<=1'b1;
29046: pixelout<=1'b1;
29047: pixelout<=1'b1;
29048: pixelout<=1'b1;
29049: pixelout<=1'b1;
29050: pixelout<=1'b1;
29051: pixelout<=1'b1;
29052: pixelout<=1'b1;
29053: pixelout<=1'b1;
29054: pixelout<=1'b1;
29055: pixelout<=1'b1;
29056: pixelout<=1'b1;
29057: pixelout<=1'b1;
29058: pixelout<=1'b1;
29059: pixelout<=1'b1;
29060: pixelout<=1'b1;
29061: pixelout<=1'b1;
29062: pixelout<=1'b1;
29063: pixelout<=1'b1;
29064: pixelout<=1'b1;
29065: pixelout<=1'b1;
29066: pixelout<=1'b1;
29067: pixelout<=1'b1;
29068: pixelout<=1'b1;
29069: pixelout<=1'b1;
29070: pixelout<=1'b1;
29071: pixelout<=1'b1;
29072: pixelout<=1'b1;
29073: pixelout<=1'b1;
29074: pixelout<=1'b1;
29075: pixelout<=1'b1;
29076: pixelout<=1'b1;
29077: pixelout<=1'b1;
29078: pixelout<=1'b1;
29079: pixelout<=1'b1;
29080: pixelout<=1'b1;
29081: pixelout<=1'b1;
29082: pixelout<=1'b1;
29083: pixelout<=1'b1;
29084: pixelout<=1'b1;
29085: pixelout<=1'b1;
29086: pixelout<=1'b1;
29087: pixelout<=1'b1;
29088: pixelout<=1'b1;
29089: pixelout<=1'b1;
29090: pixelout<=1'b1;
29091: pixelout<=1'b1;
29092: pixelout<=1'b1;
29093: pixelout<=1'b1;
29094: pixelout<=1'b1;
29095: pixelout<=1'b1;
29096: pixelout<=1'b1;
29097: pixelout<=1'b1;
29098: pixelout<=1'b1;
29099: pixelout<=1'b1;
29100: pixelout<=1'b1;
29101: pixelout<=1'b1;
29102: pixelout<=1'b1;
29103: pixelout<=1'b1;
29104: pixelout<=1'b1;
29105: pixelout<=1'b1;
29106: pixelout<=1'b1;
29107: pixelout<=1'b1;
29108: pixelout<=1'b1;
29109: pixelout<=1'b1;
29110: pixelout<=1'b1;
29111: pixelout<=1'b1;
29112: pixelout<=1'b1;
29113: pixelout<=1'b1;
29114: pixelout<=1'b1;
29115: pixelout<=1'b1;
29116: pixelout<=1'b1;
29117: pixelout<=1'b1;
29118: pixelout<=1'b1;
29119: pixelout<=1'b1;
29120: pixelout<=1'b1;
29121: pixelout<=1'b1;
29122: pixelout<=1'b1;
29123: pixelout<=1'b1;
29124: pixelout<=1'b1;
29125: pixelout<=1'b1;
29126: pixelout<=1'b1;
29127: pixelout<=1'b1;
29128: pixelout<=1'b1;
29129: pixelout<=1'b1;
29130: pixelout<=1'b1;
29131: pixelout<=1'b1;
29132: pixelout<=1'b1;
29133: pixelout<=1'b1;
29134: pixelout<=1'b1;
29135: pixelout<=1'b1;
29136: pixelout<=1'b1;
29137: pixelout<=1'b1;
29138: pixelout<=1'b1;
29139: pixelout<=1'b1;
29140: pixelout<=1'b1;
29141: pixelout<=1'b1;
29142: pixelout<=1'b1;
29143: pixelout<=1'b1;
29144: pixelout<=1'b1;
29145: pixelout<=1'b1;
29146: pixelout<=1'b1;
29147: pixelout<=1'b1;
29148: pixelout<=1'b1;
29149: pixelout<=1'b1;
29150: pixelout<=1'b1;
29151: pixelout<=1'b1;
29152: pixelout<=1'b1;
29153: pixelout<=1'b1;
29154: pixelout<=1'b1;
29155: pixelout<=1'b1;
29156: pixelout<=1'b1;
29157: pixelout<=1'b1;
29158: pixelout<=1'b1;
29159: pixelout<=1'b1;
29160: pixelout<=1'b1;
29161: pixelout<=1'b1;
29162: pixelout<=1'b1;
29163: pixelout<=1'b1;
29164: pixelout<=1'b1;
29165: pixelout<=1'b1;
29166: pixelout<=1'b1;
29167: pixelout<=1'b1;
29168: pixelout<=1'b1;
29169: pixelout<=1'b1;
29170: pixelout<=1'b1;
29171: pixelout<=1'b1;
29172: pixelout<=1'b1;
29173: pixelout<=1'b1;
29174: pixelout<=1'b1;
29175: pixelout<=1'b1;
29176: pixelout<=1'b1;
29177: pixelout<=1'b1;
29178: pixelout<=1'b1;
29179: pixelout<=1'b1;
29180: pixelout<=1'b1;
29181: pixelout<=1'b1;
29182: pixelout<=1'b1;
29183: pixelout<=1'b1;
29184: pixelout<=1'b1;
29185: pixelout<=1'b1;
29186: pixelout<=1'b1;
29187: pixelout<=1'b1;
29188: pixelout<=1'b1;
29189: pixelout<=1'b1;
29190: pixelout<=1'b1;
29191: pixelout<=1'b1;
29192: pixelout<=1'b1;
29193: pixelout<=1'b1;
29194: pixelout<=1'b1;
29195: pixelout<=1'b1;
29196: pixelout<=1'b1;
29197: pixelout<=1'b1;
29198: pixelout<=1'b1;
29199: pixelout<=1'b1;
29200: pixelout<=1'b1;
29201: pixelout<=1'b1;
29202: pixelout<=1'b1;
29203: pixelout<=1'b1;
29204: pixelout<=1'b1;
29205: pixelout<=1'b1;
29206: pixelout<=1'b1;
29207: pixelout<=1'b1;
29208: pixelout<=1'b1;
29209: pixelout<=1'b1;
29210: pixelout<=1'b1;
29211: pixelout<=1'b1;
29212: pixelout<=1'b1;
29213: pixelout<=1'b1;
29214: pixelout<=1'b1;
29215: pixelout<=1'b1;
29216: pixelout<=1'b1;
29217: pixelout<=1'b1;
29218: pixelout<=1'b1;
29219: pixelout<=1'b1;
29220: pixelout<=1'b1;
29221: pixelout<=1'b1;
29222: pixelout<=1'b1;
29223: pixelout<=1'b1;
29224: pixelout<=1'b1;
29225: pixelout<=1'b1;
29226: pixelout<=1'b1;
29227: pixelout<=1'b1;
29228: pixelout<=1'b1;
29229: pixelout<=1'b1;
29230: pixelout<=1'b1;
29231: pixelout<=1'b1;
29232: pixelout<=1'b1;
29233: pixelout<=1'b1;
29234: pixelout<=1'b1;
29235: pixelout<=1'b1;
29236: pixelout<=1'b1;
29237: pixelout<=1'b1;
29238: pixelout<=1'b1;
29239: pixelout<=1'b1;
29240: pixelout<=1'b1;
29241: pixelout<=1'b1;
29242: pixelout<=1'b1;
29243: pixelout<=1'b1;
29244: pixelout<=1'b1;
29245: pixelout<=1'b1;
29246: pixelout<=1'b1;
29247: pixelout<=1'b1;
29248: pixelout<=1'b1;
29249: pixelout<=1'b1;
29250: pixelout<=1'b1;
29251: pixelout<=1'b1;
29252: pixelout<=1'b1;
29253: pixelout<=1'b1;
29254: pixelout<=1'b1;
29255: pixelout<=1'b1;
29256: pixelout<=1'b1;
29257: pixelout<=1'b1;
29258: pixelout<=1'b1;
29259: pixelout<=1'b1;
29260: pixelout<=1'b1;
29261: pixelout<=1'b1;
29262: pixelout<=1'b1;
29263: pixelout<=1'b1;
29264: pixelout<=1'b1;
29265: pixelout<=1'b1;
29266: pixelout<=1'b1;
29267: pixelout<=1'b1;
29268: pixelout<=1'b1;
29269: pixelout<=1'b1;
29270: pixelout<=1'b1;
29271: pixelout<=1'b1;
29272: pixelout<=1'b1;
29273: pixelout<=1'b1;
29274: pixelout<=1'b1;
29275: pixelout<=1'b1;
29276: pixelout<=1'b1;
29277: pixelout<=1'b1;
29278: pixelout<=1'b1;
29279: pixelout<=1'b1;
29280: pixelout<=1'b1;
29281: pixelout<=1'b1;
29282: pixelout<=1'b1;
29283: pixelout<=1'b1;
29284: pixelout<=1'b1;
29285: pixelout<=1'b1;
29286: pixelout<=1'b1;
29287: pixelout<=1'b1;
29288: pixelout<=1'b1;
29289: pixelout<=1'b1;
29290: pixelout<=1'b1;
29291: pixelout<=1'b1;
29292: pixelout<=1'b1;
29293: pixelout<=1'b1;
29294: pixelout<=1'b1;
29295: pixelout<=1'b1;
29296: pixelout<=1'b1;
29297: pixelout<=1'b1;
29298: pixelout<=1'b1;
29299: pixelout<=1'b1;
29300: pixelout<=1'b1;
29301: pixelout<=1'b1;
29302: pixelout<=1'b1;
29303: pixelout<=1'b1;
29304: pixelout<=1'b1;
29305: pixelout<=1'b1;
29306: pixelout<=1'b1;
29307: pixelout<=1'b1;
29308: pixelout<=1'b1;
29309: pixelout<=1'b1;
29310: pixelout<=1'b1;
29311: pixelout<=1'b1;
29312: pixelout<=1'b1;
29313: pixelout<=1'b1;
29314: pixelout<=1'b1;
29315: pixelout<=1'b1;
29316: pixelout<=1'b1;
29317: pixelout<=1'b1;
29318: pixelout<=1'b1;
29319: pixelout<=1'b1;
29320: pixelout<=1'b1;
29321: pixelout<=1'b1;
29322: pixelout<=1'b1;
29323: pixelout<=1'b1;
29324: pixelout<=1'b1;
29325: pixelout<=1'b1;
29326: pixelout<=1'b1;
29327: pixelout<=1'b1;
29328: pixelout<=1'b1;
29329: pixelout<=1'b1;
29330: pixelout<=1'b1;
29331: pixelout<=1'b1;
29332: pixelout<=1'b1;
29333: pixelout<=1'b1;
29334: pixelout<=1'b1;
29335: pixelout<=1'b1;
29336: pixelout<=1'b1;
29337: pixelout<=1'b1;
29338: pixelout<=1'b1;
29339: pixelout<=1'b1;
29340: pixelout<=1'b1;
29341: pixelout<=1'b1;
29342: pixelout<=1'b1;
29343: pixelout<=1'b1;
29344: pixelout<=1'b1;
29345: pixelout<=1'b1;
29346: pixelout<=1'b1;
29347: pixelout<=1'b1;
29348: pixelout<=1'b1;
29349: pixelout<=1'b1;
29350: pixelout<=1'b1;
29351: pixelout<=1'b1;
29352: pixelout<=1'b1;
29353: pixelout<=1'b1;
29354: pixelout<=1'b1;
29355: pixelout<=1'b1;
29356: pixelout<=1'b1;
29357: pixelout<=1'b1;
29358: pixelout<=1'b1;
29359: pixelout<=1'b1;
29360: pixelout<=1'b1;
29361: pixelout<=1'b1;
29362: pixelout<=1'b1;
29363: pixelout<=1'b1;
29364: pixelout<=1'b1;
29365: pixelout<=1'b1;
29366: pixelout<=1'b1;
29367: pixelout<=1'b1;
29368: pixelout<=1'b1;
29369: pixelout<=1'b1;
29370: pixelout<=1'b1;
29371: pixelout<=1'b1;
29372: pixelout<=1'b1;
29373: pixelout<=1'b1;
29374: pixelout<=1'b1;
29375: pixelout<=1'b1;
29376: pixelout<=1'b1;
29377: pixelout<=1'b1;
29378: pixelout<=1'b1;
29379: pixelout<=1'b1;
29380: pixelout<=1'b1;
29381: pixelout<=1'b1;
29382: pixelout<=1'b1;
29383: pixelout<=1'b1;
29384: pixelout<=1'b1;
29385: pixelout<=1'b1;
29386: pixelout<=1'b1;
29387: pixelout<=1'b1;
29388: pixelout<=1'b1;
29389: pixelout<=1'b1;
29390: pixelout<=1'b1;
29391: pixelout<=1'b1;
29392: pixelout<=1'b1;
29393: pixelout<=1'b1;
29394: pixelout<=1'b1;
29395: pixelout<=1'b1;
29396: pixelout<=1'b1;
29397: pixelout<=1'b1;
29398: pixelout<=1'b1;
29399: pixelout<=1'b1;
29400: pixelout<=1'b1;
29401: pixelout<=1'b1;
29402: pixelout<=1'b1;
29403: pixelout<=1'b1;
29404: pixelout<=1'b1;
29405: pixelout<=1'b1;
29406: pixelout<=1'b1;
29407: pixelout<=1'b1;
29408: pixelout<=1'b1;
29409: pixelout<=1'b1;
29410: pixelout<=1'b1;
29411: pixelout<=1'b1;
29412: pixelout<=1'b1;
29413: pixelout<=1'b1;
29414: pixelout<=1'b1;
29415: pixelout<=1'b1;
29416: pixelout<=1'b1;
29417: pixelout<=1'b1;
29418: pixelout<=1'b1;
29419: pixelout<=1'b1;
29420: pixelout<=1'b1;
29421: pixelout<=1'b1;
29422: pixelout<=1'b1;
29423: pixelout<=1'b1;
29424: pixelout<=1'b1;
29425: pixelout<=1'b1;
29426: pixelout<=1'b1;
29427: pixelout<=1'b1;
29428: pixelout<=1'b1;
29429: pixelout<=1'b1;
29430: pixelout<=1'b1;
29431: pixelout<=1'b1;
29432: pixelout<=1'b1;
29433: pixelout<=1'b1;
29434: pixelout<=1'b1;
29435: pixelout<=1'b1;
29436: pixelout<=1'b1;
29437: pixelout<=1'b1;
29438: pixelout<=1'b1;
29439: pixelout<=1'b1;
29440: pixelout<=1'b1;
29441: pixelout<=1'b1;
29442: pixelout<=1'b1;
29443: pixelout<=1'b1;
29444: pixelout<=1'b1;
29445: pixelout<=1'b1;
29446: pixelout<=1'b1;
29447: pixelout<=1'b1;
29448: pixelout<=1'b1;
29449: pixelout<=1'b1;
29450: pixelout<=1'b1;
29451: pixelout<=1'b1;
29452: pixelout<=1'b1;
29453: pixelout<=1'b1;
29454: pixelout<=1'b1;
29455: pixelout<=1'b1;
29456: pixelout<=1'b1;
29457: pixelout<=1'b1;
29458: pixelout<=1'b1;
29459: pixelout<=1'b1;
29460: pixelout<=1'b1;
29461: pixelout<=1'b1;
29462: pixelout<=1'b1;
29463: pixelout<=1'b1;
29464: pixelout<=1'b1;
29465: pixelout<=1'b1;
29466: pixelout<=1'b1;
29467: pixelout<=1'b1;
29468: pixelout<=1'b1;
29469: pixelout<=1'b1;
29470: pixelout<=1'b1;
29471: pixelout<=1'b1;
29472: pixelout<=1'b1;
29473: pixelout<=1'b1;
29474: pixelout<=1'b1;
29475: pixelout<=1'b1;
29476: pixelout<=1'b1;
29477: pixelout<=1'b1;
29478: pixelout<=1'b1;
29479: pixelout<=1'b1;
29480: pixelout<=1'b1;
29481: pixelout<=1'b1;
29482: pixelout<=1'b1;
29483: pixelout<=1'b1;
29484: pixelout<=1'b1;
29485: pixelout<=1'b1;
29486: pixelout<=1'b1;
29487: pixelout<=1'b1;
29488: pixelout<=1'b1;
29489: pixelout<=1'b1;
29490: pixelout<=1'b1;
29491: pixelout<=1'b1;
29492: pixelout<=1'b1;
29493: pixelout<=1'b1;
29494: pixelout<=1'b1;
29495: pixelout<=1'b1;
29496: pixelout<=1'b1;
29497: pixelout<=1'b1;
29498: pixelout<=1'b1;
29499: pixelout<=1'b1;
29500: pixelout<=1'b1;
29501: pixelout<=1'b1;
29502: pixelout<=1'b1;
29503: pixelout<=1'b1;
29504: pixelout<=1'b1;
29505: pixelout<=1'b1;
29506: pixelout<=1'b1;
29507: pixelout<=1'b1;
29508: pixelout<=1'b1;
29509: pixelout<=1'b1;
29510: pixelout<=1'b1;
29511: pixelout<=1'b1;
29512: pixelout<=1'b1;
29513: pixelout<=1'b1;
29514: pixelout<=1'b1;
29515: pixelout<=1'b1;
29516: pixelout<=1'b1;
29517: pixelout<=1'b1;
29518: pixelout<=1'b1;
29519: pixelout<=1'b1;
29520: pixelout<=1'b1;
29521: pixelout<=1'b1;
29522: pixelout<=1'b1;
29523: pixelout<=1'b1;
29524: pixelout<=1'b1;
29525: pixelout<=1'b1;
29526: pixelout<=1'b1;
29527: pixelout<=1'b1;
29528: pixelout<=1'b1;
29529: pixelout<=1'b1;
29530: pixelout<=1'b1;
29531: pixelout<=1'b1;
29532: pixelout<=1'b1;
29533: pixelout<=1'b1;
29534: pixelout<=1'b1;
29535: pixelout<=1'b1;
29536: pixelout<=1'b1;
29537: pixelout<=1'b1;
29538: pixelout<=1'b1;
29539: pixelout<=1'b1;
29540: pixelout<=1'b1;
29541: pixelout<=1'b1;
29542: pixelout<=1'b1;
29543: pixelout<=1'b1;
29544: pixelout<=1'b1;
29545: pixelout<=1'b1;
29546: pixelout<=1'b1;
29547: pixelout<=1'b1;
29548: pixelout<=1'b1;
29549: pixelout<=1'b1;
29550: pixelout<=1'b1;
29551: pixelout<=1'b1;
29552: pixelout<=1'b1;
29553: pixelout<=1'b1;
29554: pixelout<=1'b1;
29555: pixelout<=1'b1;
29556: pixelout<=1'b1;
29557: pixelout<=1'b1;
29558: pixelout<=1'b1;
29559: pixelout<=1'b1;
29560: pixelout<=1'b1;
29561: pixelout<=1'b1;
29562: pixelout<=1'b1;
29563: pixelout<=1'b1;
29564: pixelout<=1'b1;
29565: pixelout<=1'b1;
29566: pixelout<=1'b1;
29567: pixelout<=1'b1;
29568: pixelout<=1'b1;
29569: pixelout<=1'b1;
29570: pixelout<=1'b1;
29571: pixelout<=1'b1;
29572: pixelout<=1'b1;
29573: pixelout<=1'b1;
29574: pixelout<=1'b1;
29575: pixelout<=1'b1;
29576: pixelout<=1'b1;
29577: pixelout<=1'b1;
29578: pixelout<=1'b1;
29579: pixelout<=1'b1;
29580: pixelout<=1'b1;
29581: pixelout<=1'b1;
29582: pixelout<=1'b1;
29583: pixelout<=1'b1;
29584: pixelout<=1'b1;
29585: pixelout<=1'b1;
29586: pixelout<=1'b1;
29587: pixelout<=1'b1;
29588: pixelout<=1'b1;
29589: pixelout<=1'b1;
29590: pixelout<=1'b1;
29591: pixelout<=1'b1;
29592: pixelout<=1'b1;
29593: pixelout<=1'b1;
29594: pixelout<=1'b1;
29595: pixelout<=1'b1;
29596: pixelout<=1'b1;
29597: pixelout<=1'b1;
29598: pixelout<=1'b1;
29599: pixelout<=1'b1;
29600: pixelout<=1'b1;
29601: pixelout<=1'b1;
29602: pixelout<=1'b1;
29603: pixelout<=1'b1;
29604: pixelout<=1'b1;
29605: pixelout<=1'b1;
29606: pixelout<=1'b1;
29607: pixelout<=1'b1;
29608: pixelout<=1'b1;
29609: pixelout<=1'b1;
29610: pixelout<=1'b1;
29611: pixelout<=1'b1;
29612: pixelout<=1'b1;
29613: pixelout<=1'b1;
29614: pixelout<=1'b1;
29615: pixelout<=1'b1;
29616: pixelout<=1'b1;
29617: pixelout<=1'b1;
29618: pixelout<=1'b1;
29619: pixelout<=1'b1;
29620: pixelout<=1'b1;
29621: pixelout<=1'b1;
29622: pixelout<=1'b1;
29623: pixelout<=1'b1;
29624: pixelout<=1'b1;
29625: pixelout<=1'b1;
29626: pixelout<=1'b1;
29627: pixelout<=1'b1;
29628: pixelout<=1'b1;
29629: pixelout<=1'b1;
29630: pixelout<=1'b1;
29631: pixelout<=1'b1;
29632: pixelout<=1'b1;
29633: pixelout<=1'b1;
29634: pixelout<=1'b1;
29635: pixelout<=1'b1;
29636: pixelout<=1'b1;
29637: pixelout<=1'b1;
29638: pixelout<=1'b1;
29639: pixelout<=1'b1;
29640: pixelout<=1'b1;
29641: pixelout<=1'b1;
29642: pixelout<=1'b1;
29643: pixelout<=1'b1;
29644: pixelout<=1'b1;
29645: pixelout<=1'b1;
29646: pixelout<=1'b1;
29647: pixelout<=1'b1;
29648: pixelout<=1'b1;
29649: pixelout<=1'b1;
29650: pixelout<=1'b1;
29651: pixelout<=1'b1;
29652: pixelout<=1'b1;
29653: pixelout<=1'b1;
29654: pixelout<=1'b1;
29655: pixelout<=1'b1;
29656: pixelout<=1'b1;
29657: pixelout<=1'b1;
29658: pixelout<=1'b1;
29659: pixelout<=1'b1;
29660: pixelout<=1'b1;
29661: pixelout<=1'b1;
29662: pixelout<=1'b1;
29663: pixelout<=1'b1;
29664: pixelout<=1'b1;
29665: pixelout<=1'b1;
29666: pixelout<=1'b1;
29667: pixelout<=1'b1;
29668: pixelout<=1'b1;
29669: pixelout<=1'b1;
29670: pixelout<=1'b1;
29671: pixelout<=1'b1;
29672: pixelout<=1'b1;
29673: pixelout<=1'b1;
29674: pixelout<=1'b1;
29675: pixelout<=1'b1;
29676: pixelout<=1'b1;
29677: pixelout<=1'b1;
29678: pixelout<=1'b1;
29679: pixelout<=1'b1;
29680: pixelout<=1'b1;
29681: pixelout<=1'b1;
29682: pixelout<=1'b1;
29683: pixelout<=1'b1;
29684: pixelout<=1'b1;
29685: pixelout<=1'b1;
29686: pixelout<=1'b1;
29687: pixelout<=1'b1;
29688: pixelout<=1'b1;
29689: pixelout<=1'b1;
29690: pixelout<=1'b1;
29691: pixelout<=1'b1;
29692: pixelout<=1'b1;
29693: pixelout<=1'b1;
29694: pixelout<=1'b1;
29695: pixelout<=1'b1;
29696: pixelout<=1'b1;
29697: pixelout<=1'b1;
29698: pixelout<=1'b1;
29699: pixelout<=1'b1;
29700: pixelout<=1'b1;
29701: pixelout<=1'b1;
29702: pixelout<=1'b1;
29703: pixelout<=1'b1;
29704: pixelout<=1'b1;
29705: pixelout<=1'b1;
29706: pixelout<=1'b1;
29707: pixelout<=1'b1;
29708: pixelout<=1'b1;
29709: pixelout<=1'b1;
29710: pixelout<=1'b1;
29711: pixelout<=1'b1;
29712: pixelout<=1'b1;
29713: pixelout<=1'b1;
29714: pixelout<=1'b1;
29715: pixelout<=1'b1;
29716: pixelout<=1'b1;
29717: pixelout<=1'b1;
29718: pixelout<=1'b1;
29719: pixelout<=1'b1;
29720: pixelout<=1'b1;
29721: pixelout<=1'b1;
29722: pixelout<=1'b1;
29723: pixelout<=1'b1;
29724: pixelout<=1'b1;
29725: pixelout<=1'b1;
29726: pixelout<=1'b1;
29727: pixelout<=1'b1;
29728: pixelout<=1'b1;
29729: pixelout<=1'b1;
29730: pixelout<=1'b1;
29731: pixelout<=1'b1;
29732: pixelout<=1'b1;
29733: pixelout<=1'b1;
29734: pixelout<=1'b1;
29735: pixelout<=1'b1;
29736: pixelout<=1'b1;
29737: pixelout<=1'b1;
29738: pixelout<=1'b1;
29739: pixelout<=1'b1;
29740: pixelout<=1'b1;
29741: pixelout<=1'b1;
29742: pixelout<=1'b1;
29743: pixelout<=1'b1;
29744: pixelout<=1'b1;
29745: pixelout<=1'b1;
29746: pixelout<=1'b1;
29747: pixelout<=1'b1;
29748: pixelout<=1'b1;
29749: pixelout<=1'b1;
29750: pixelout<=1'b1;
29751: pixelout<=1'b1;
29752: pixelout<=1'b1;
29753: pixelout<=1'b1;
29754: pixelout<=1'b1;
29755: pixelout<=1'b1;
29756: pixelout<=1'b1;
29757: pixelout<=1'b1;
29758: pixelout<=1'b1;
29759: pixelout<=1'b1;
29760: pixelout<=1'b1;
29761: pixelout<=1'b1;
29762: pixelout<=1'b1;
29763: pixelout<=1'b1;
29764: pixelout<=1'b1;
29765: pixelout<=1'b1;
29766: pixelout<=1'b1;
29767: pixelout<=1'b1;
29768: pixelout<=1'b1;
29769: pixelout<=1'b1;
29770: pixelout<=1'b1;
29771: pixelout<=1'b1;
29772: pixelout<=1'b1;
29773: pixelout<=1'b1;
29774: pixelout<=1'b1;
29775: pixelout<=1'b1;
29776: pixelout<=1'b1;
29777: pixelout<=1'b1;
29778: pixelout<=1'b1;
29779: pixelout<=1'b1;
29780: pixelout<=1'b1;
29781: pixelout<=1'b1;
29782: pixelout<=1'b1;
29783: pixelout<=1'b1;
29784: pixelout<=1'b1;
29785: pixelout<=1'b1;
29786: pixelout<=1'b1;
29787: pixelout<=1'b1;
29788: pixelout<=1'b1;
29789: pixelout<=1'b1;
29790: pixelout<=1'b1;
29791: pixelout<=1'b1;
29792: pixelout<=1'b1;
29793: pixelout<=1'b1;
29794: pixelout<=1'b1;
29795: pixelout<=1'b1;
29796: pixelout<=1'b1;
29797: pixelout<=1'b1;
29798: pixelout<=1'b1;
29799: pixelout<=1'b1;
29800: pixelout<=1'b1;
29801: pixelout<=1'b1;
29802: pixelout<=1'b1;
29803: pixelout<=1'b1;
29804: pixelout<=1'b1;
29805: pixelout<=1'b1;
29806: pixelout<=1'b1;
29807: pixelout<=1'b1;
29808: pixelout<=1'b1;
29809: pixelout<=1'b1;
29810: pixelout<=1'b1;
29811: pixelout<=1'b1;
29812: pixelout<=1'b1;
29813: pixelout<=1'b1;
29814: pixelout<=1'b1;
29815: pixelout<=1'b1;
29816: pixelout<=1'b1;
29817: pixelout<=1'b1;
29818: pixelout<=1'b1;
29819: pixelout<=1'b1;
29820: pixelout<=1'b1;
29821: pixelout<=1'b1;
29822: pixelout<=1'b1;
29823: pixelout<=1'b1;
29824: pixelout<=1'b1;
29825: pixelout<=1'b1;
29826: pixelout<=1'b1;
29827: pixelout<=1'b1;
29828: pixelout<=1'b1;
29829: pixelout<=1'b1;
29830: pixelout<=1'b1;
29831: pixelout<=1'b1;
29832: pixelout<=1'b1;
29833: pixelout<=1'b1;
29834: pixelout<=1'b1;
29835: pixelout<=1'b1;
29836: pixelout<=1'b1;
29837: pixelout<=1'b1;
29838: pixelout<=1'b1;
29839: pixelout<=1'b1;
29840: pixelout<=1'b1;
29841: pixelout<=1'b1;
29842: pixelout<=1'b1;
29843: pixelout<=1'b1;
29844: pixelout<=1'b1;
29845: pixelout<=1'b1;
29846: pixelout<=1'b1;
29847: pixelout<=1'b1;
29848: pixelout<=1'b1;
29849: pixelout<=1'b1;
29850: pixelout<=1'b1;
29851: pixelout<=1'b1;
29852: pixelout<=1'b1;
29853: pixelout<=1'b1;
29854: pixelout<=1'b1;
29855: pixelout<=1'b1;
29856: pixelout<=1'b1;
29857: pixelout<=1'b1;
29858: pixelout<=1'b1;
29859: pixelout<=1'b1;
29860: pixelout<=1'b1;
29861: pixelout<=1'b1;
29862: pixelout<=1'b1;
29863: pixelout<=1'b1;
29864: pixelout<=1'b1;
29865: pixelout<=1'b1;
29866: pixelout<=1'b1;
29867: pixelout<=1'b1;
29868: pixelout<=1'b1;
29869: pixelout<=1'b1;
29870: pixelout<=1'b1;
29871: pixelout<=1'b1;
29872: pixelout<=1'b1;
29873: pixelout<=1'b1;
29874: pixelout<=1'b1;
29875: pixelout<=1'b1;
29876: pixelout<=1'b1;
29877: pixelout<=1'b1;
29878: pixelout<=1'b1;
29879: pixelout<=1'b1;
29880: pixelout<=1'b1;
29881: pixelout<=1'b1;
29882: pixelout<=1'b1;
29883: pixelout<=1'b1;
29884: pixelout<=1'b1;
29885: pixelout<=1'b1;
29886: pixelout<=1'b1;
29887: pixelout<=1'b1;
29888: pixelout<=1'b1;
29889: pixelout<=1'b1;
29890: pixelout<=1'b1;
29891: pixelout<=1'b1;
29892: pixelout<=1'b1;
29893: pixelout<=1'b1;
29894: pixelout<=1'b1;
29895: pixelout<=1'b1;
29896: pixelout<=1'b1;
29897: pixelout<=1'b1;
29898: pixelout<=1'b1;
29899: pixelout<=1'b1;
29900: pixelout<=1'b1;
29901: pixelout<=1'b1;
29902: pixelout<=1'b1;
29903: pixelout<=1'b1;
29904: pixelout<=1'b1;
29905: pixelout<=1'b1;
29906: pixelout<=1'b1;
29907: pixelout<=1'b1;
29908: pixelout<=1'b1;
29909: pixelout<=1'b1;
29910: pixelout<=1'b1;
29911: pixelout<=1'b1;
29912: pixelout<=1'b1;
29913: pixelout<=1'b1;
29914: pixelout<=1'b1;
29915: pixelout<=1'b1;
29916: pixelout<=1'b1;
29917: pixelout<=1'b1;
29918: pixelout<=1'b1;
29919: pixelout<=1'b1;
29920: pixelout<=1'b1;
29921: pixelout<=1'b1;
29922: pixelout<=1'b1;
29923: pixelout<=1'b1;
29924: pixelout<=1'b1;
29925: pixelout<=1'b1;
29926: pixelout<=1'b1;
29927: pixelout<=1'b1;
29928: pixelout<=1'b1;
29929: pixelout<=1'b1;
29930: pixelout<=1'b1;
29931: pixelout<=1'b1;
29932: pixelout<=1'b1;
29933: pixelout<=1'b1;
29934: pixelout<=1'b1;
29935: pixelout<=1'b1;
29936: pixelout<=1'b1;
29937: pixelout<=1'b1;
29938: pixelout<=1'b1;
29939: pixelout<=1'b1;
29940: pixelout<=1'b1;
29941: pixelout<=1'b1;
29942: pixelout<=1'b1;
29943: pixelout<=1'b1;
29944: pixelout<=1'b1;
29945: pixelout<=1'b1;
29946: pixelout<=1'b1;
29947: pixelout<=1'b1;
29948: pixelout<=1'b1;
29949: pixelout<=1'b1;
29950: pixelout<=1'b1;
29951: pixelout<=1'b1;
29952: pixelout<=1'b1;
29953: pixelout<=1'b1;
29954: pixelout<=1'b1;
29955: pixelout<=1'b1;
29956: pixelout<=1'b1;
29957: pixelout<=1'b1;
29958: pixelout<=1'b1;
29959: pixelout<=1'b1;
29960: pixelout<=1'b1;
29961: pixelout<=1'b1;
29962: pixelout<=1'b1;
29963: pixelout<=1'b1;
29964: pixelout<=1'b1;
29965: pixelout<=1'b1;
29966: pixelout<=1'b1;
29967: pixelout<=1'b1;
29968: pixelout<=1'b1;
29969: pixelout<=1'b1;
29970: pixelout<=1'b1;
29971: pixelout<=1'b1;
29972: pixelout<=1'b1;
29973: pixelout<=1'b1;
29974: pixelout<=1'b1;
29975: pixelout<=1'b1;
29976: pixelout<=1'b1;
29977: pixelout<=1'b1;
29978: pixelout<=1'b1;
29979: pixelout<=1'b1;
29980: pixelout<=1'b1;
29981: pixelout<=1'b1;
29982: pixelout<=1'b1;
29983: pixelout<=1'b1;
29984: pixelout<=1'b1;
29985: pixelout<=1'b1;
29986: pixelout<=1'b1;
29987: pixelout<=1'b1;
29988: pixelout<=1'b1;
29989: pixelout<=1'b1;
29990: pixelout<=1'b1;
29991: pixelout<=1'b1;
29992: pixelout<=1'b1;
29993: pixelout<=1'b1;
29994: pixelout<=1'b1;
29995: pixelout<=1'b1;
29996: pixelout<=1'b1;
29997: pixelout<=1'b1;
29998: pixelout<=1'b1;
29999: pixelout<=1'b1;
30000: pixelout<=1'b1;
30001: pixelout<=1'b1;
30002: pixelout<=1'b1;
30003: pixelout<=1'b1;
30004: pixelout<=1'b1;
30005: pixelout<=1'b1;
30006: pixelout<=1'b1;
30007: pixelout<=1'b1;
30008: pixelout<=1'b1;
30009: pixelout<=1'b1;
30010: pixelout<=1'b1;
30011: pixelout<=1'b1;
30012: pixelout<=1'b1;
30013: pixelout<=1'b1;
30014: pixelout<=1'b1;
30015: pixelout<=1'b1;
30016: pixelout<=1'b1;
30017: pixelout<=1'b1;
30018: pixelout<=1'b1;
30019: pixelout<=1'b1;
30020: pixelout<=1'b1;
30021: pixelout<=1'b1;
30022: pixelout<=1'b1;
30023: pixelout<=1'b1;
30024: pixelout<=1'b1;
30025: pixelout<=1'b1;
30026: pixelout<=1'b1;
30027: pixelout<=1'b1;
30028: pixelout<=1'b1;
30029: pixelout<=1'b1;
30030: pixelout<=1'b1;
30031: pixelout<=1'b1;
30032: pixelout<=1'b1;
30033: pixelout<=1'b1;
30034: pixelout<=1'b1;
30035: pixelout<=1'b1;
30036: pixelout<=1'b1;
30037: pixelout<=1'b1;
30038: pixelout<=1'b1;
30039: pixelout<=1'b1;
30040: pixelout<=1'b1;
30041: pixelout<=1'b1;
30042: pixelout<=1'b1;
30043: pixelout<=1'b1;
30044: pixelout<=1'b1;
30045: pixelout<=1'b1;
30046: pixelout<=1'b1;
30047: pixelout<=1'b1;
30048: pixelout<=1'b1;
30049: pixelout<=1'b1;
30050: pixelout<=1'b1;
30051: pixelout<=1'b1;
30052: pixelout<=1'b1;
30053: pixelout<=1'b1;
30054: pixelout<=1'b1;
30055: pixelout<=1'b1;
30056: pixelout<=1'b1;
30057: pixelout<=1'b1;
30058: pixelout<=1'b1;
30059: pixelout<=1'b1;
30060: pixelout<=1'b1;
30061: pixelout<=1'b1;
30062: pixelout<=1'b1;
30063: pixelout<=1'b1;
30064: pixelout<=1'b1;
30065: pixelout<=1'b1;
30066: pixelout<=1'b1;
30067: pixelout<=1'b1;
30068: pixelout<=1'b1;
30069: pixelout<=1'b1;
30070: pixelout<=1'b1;
30071: pixelout<=1'b1;
30072: pixelout<=1'b1;
30073: pixelout<=1'b1;
30074: pixelout<=1'b1;
30075: pixelout<=1'b1;
30076: pixelout<=1'b1;
30077: pixelout<=1'b1;
30078: pixelout<=1'b1;
30079: pixelout<=1'b1;
30080: pixelout<=1'b1;
30081: pixelout<=1'b1;
30082: pixelout<=1'b1;
30083: pixelout<=1'b1;
30084: pixelout<=1'b1;
30085: pixelout<=1'b1;
30086: pixelout<=1'b1;
30087: pixelout<=1'b1;
30088: pixelout<=1'b1;
30089: pixelout<=1'b1;
30090: pixelout<=1'b1;
30091: pixelout<=1'b1;
30092: pixelout<=1'b1;
30093: pixelout<=1'b1;
30094: pixelout<=1'b1;
30095: pixelout<=1'b1;
30096: pixelout<=1'b1;
30097: pixelout<=1'b1;
30098: pixelout<=1'b1;
30099: pixelout<=1'b1;
30100: pixelout<=1'b1;
30101: pixelout<=1'b1;
30102: pixelout<=1'b1;
30103: pixelout<=1'b1;
30104: pixelout<=1'b1;
30105: pixelout<=1'b1;
30106: pixelout<=1'b1;
30107: pixelout<=1'b1;
30108: pixelout<=1'b1;
30109: pixelout<=1'b1;
30110: pixelout<=1'b1;
30111: pixelout<=1'b1;
30112: pixelout<=1'b1;
30113: pixelout<=1'b1;
30114: pixelout<=1'b1;
30115: pixelout<=1'b1;
30116: pixelout<=1'b1;
30117: pixelout<=1'b1;
30118: pixelout<=1'b1;
30119: pixelout<=1'b1;
30120: pixelout<=1'b1;
30121: pixelout<=1'b1;
30122: pixelout<=1'b1;
30123: pixelout<=1'b1;
30124: pixelout<=1'b1;
30125: pixelout<=1'b1;
30126: pixelout<=1'b1;
30127: pixelout<=1'b1;
30128: pixelout<=1'b1;
30129: pixelout<=1'b1;
30130: pixelout<=1'b1;
30131: pixelout<=1'b1;
30132: pixelout<=1'b1;
30133: pixelout<=1'b1;
30134: pixelout<=1'b1;
30135: pixelout<=1'b1;
30136: pixelout<=1'b1;
30137: pixelout<=1'b1;
30138: pixelout<=1'b1;
30139: pixelout<=1'b1;
30140: pixelout<=1'b1;
30141: pixelout<=1'b1;
30142: pixelout<=1'b1;
30143: pixelout<=1'b1;
30144: pixelout<=1'b1;
30145: pixelout<=1'b1;
30146: pixelout<=1'b1;
30147: pixelout<=1'b1;
30148: pixelout<=1'b1;
30149: pixelout<=1'b1;
30150: pixelout<=1'b1;
30151: pixelout<=1'b1;
30152: pixelout<=1'b1;
30153: pixelout<=1'b1;
30154: pixelout<=1'b1;
30155: pixelout<=1'b1;
30156: pixelout<=1'b1;
30157: pixelout<=1'b1;
30158: pixelout<=1'b1;
30159: pixelout<=1'b1;
30160: pixelout<=1'b1;
30161: pixelout<=1'b1;
30162: pixelout<=1'b1;
30163: pixelout<=1'b1;
30164: pixelout<=1'b1;
30165: pixelout<=1'b1;
30166: pixelout<=1'b1;
30167: pixelout<=1'b1;
30168: pixelout<=1'b1;
30169: pixelout<=1'b1;
30170: pixelout<=1'b1;
30171: pixelout<=1'b1;
30172: pixelout<=1'b1;
30173: pixelout<=1'b1;
30174: pixelout<=1'b1;
30175: pixelout<=1'b1;
30176: pixelout<=1'b1;
30177: pixelout<=1'b1;
30178: pixelout<=1'b1;
30179: pixelout<=1'b1;
30180: pixelout<=1'b1;
30181: pixelout<=1'b1;
30182: pixelout<=1'b1;
30183: pixelout<=1'b1;
30184: pixelout<=1'b1;
30185: pixelout<=1'b1;
30186: pixelout<=1'b1;
30187: pixelout<=1'b1;
30188: pixelout<=1'b1;
30189: pixelout<=1'b1;
30190: pixelout<=1'b1;
30191: pixelout<=1'b1;
30192: pixelout<=1'b1;
30193: pixelout<=1'b1;
30194: pixelout<=1'b1;
30195: pixelout<=1'b1;
30196: pixelout<=1'b1;
30197: pixelout<=1'b1;
30198: pixelout<=1'b1;
30199: pixelout<=1'b1;
30200: pixelout<=1'b1;
30201: pixelout<=1'b1;
30202: pixelout<=1'b1;
30203: pixelout<=1'b1;
30204: pixelout<=1'b1;
30205: pixelout<=1'b1;
30206: pixelout<=1'b1;
30207: pixelout<=1'b1;
30208: pixelout<=1'b1;
30209: pixelout<=1'b1;
30210: pixelout<=1'b1;
30211: pixelout<=1'b1;
30212: pixelout<=1'b1;
30213: pixelout<=1'b1;
30214: pixelout<=1'b1;
30215: pixelout<=1'b1;
30216: pixelout<=1'b1;
30217: pixelout<=1'b1;
30218: pixelout<=1'b1;
30219: pixelout<=1'b1;
30220: pixelout<=1'b1;
30221: pixelout<=1'b1;
30222: pixelout<=1'b1;
30223: pixelout<=1'b1;
30224: pixelout<=1'b1;
30225: pixelout<=1'b1;
30226: pixelout<=1'b1;
30227: pixelout<=1'b1;
30228: pixelout<=1'b1;
30229: pixelout<=1'b1;
30230: pixelout<=1'b1;
30231: pixelout<=1'b1;
30232: pixelout<=1'b1;
30233: pixelout<=1'b1;
30234: pixelout<=1'b1;
30235: pixelout<=1'b1;
30236: pixelout<=1'b1;
30237: pixelout<=1'b1;
30238: pixelout<=1'b1;
30239: pixelout<=1'b1;
30240: pixelout<=1'b1;
30241: pixelout<=1'b1;
30242: pixelout<=1'b1;
30243: pixelout<=1'b1;
30244: pixelout<=1'b1;
30245: pixelout<=1'b1;
30246: pixelout<=1'b1;
30247: pixelout<=1'b1;
30248: pixelout<=1'b1;
30249: pixelout<=1'b1;
30250: pixelout<=1'b1;
30251: pixelout<=1'b1;
30252: pixelout<=1'b1;
30253: pixelout<=1'b1;
30254: pixelout<=1'b1;
30255: pixelout<=1'b1;
30256: pixelout<=1'b1;
30257: pixelout<=1'b1;
30258: pixelout<=1'b1;
30259: pixelout<=1'b1;
30260: pixelout<=1'b1;
30261: pixelout<=1'b1;
30262: pixelout<=1'b1;
30263: pixelout<=1'b1;
30264: pixelout<=1'b1;
30265: pixelout<=1'b1;
30266: pixelout<=1'b1;
30267: pixelout<=1'b1;
30268: pixelout<=1'b1;
30269: pixelout<=1'b1;
30270: pixelout<=1'b1;
30271: pixelout<=1'b1;
30272: pixelout<=1'b1;
30273: pixelout<=1'b1;
30274: pixelout<=1'b1;
30275: pixelout<=1'b1;
30276: pixelout<=1'b1;
30277: pixelout<=1'b1;
30278: pixelout<=1'b1;
30279: pixelout<=1'b1;
30280: pixelout<=1'b1;
30281: pixelout<=1'b1;
30282: pixelout<=1'b1;
30283: pixelout<=1'b1;
30284: pixelout<=1'b1;
30285: pixelout<=1'b1;
30286: pixelout<=1'b1;
30287: pixelout<=1'b1;
30288: pixelout<=1'b1;
30289: pixelout<=1'b1;
30290: pixelout<=1'b1;
30291: pixelout<=1'b1;
30292: pixelout<=1'b1;
30293: pixelout<=1'b1;
30294: pixelout<=1'b1;
30295: pixelout<=1'b1;
30296: pixelout<=1'b1;
30297: pixelout<=1'b1;
30298: pixelout<=1'b1;
30299: pixelout<=1'b1;
30300: pixelout<=1'b1;
30301: pixelout<=1'b1;
30302: pixelout<=1'b1;
30303: pixelout<=1'b1;
30304: pixelout<=1'b1;
30305: pixelout<=1'b1;
30306: pixelout<=1'b1;
30307: pixelout<=1'b1;
30308: pixelout<=1'b1;
30309: pixelout<=1'b1;
30310: pixelout<=1'b1;
30311: pixelout<=1'b1;
30312: pixelout<=1'b1;
30313: pixelout<=1'b1;
30314: pixelout<=1'b1;
30315: pixelout<=1'b1;
30316: pixelout<=1'b1;
30317: pixelout<=1'b1;
30318: pixelout<=1'b1;
30319: pixelout<=1'b1;
30320: pixelout<=1'b1;
30321: pixelout<=1'b1;
30322: pixelout<=1'b1;
30323: pixelout<=1'b1;
30324: pixelout<=1'b1;
30325: pixelout<=1'b1;
30326: pixelout<=1'b1;
30327: pixelout<=1'b1;
30328: pixelout<=1'b1;
30329: pixelout<=1'b1;
30330: pixelout<=1'b1;
30331: pixelout<=1'b1;
30332: pixelout<=1'b1;
30333: pixelout<=1'b1;
30334: pixelout<=1'b1;
30335: pixelout<=1'b1;
30336: pixelout<=1'b1;
30337: pixelout<=1'b1;
30338: pixelout<=1'b1;
30339: pixelout<=1'b1;
30340: pixelout<=1'b1;
30341: pixelout<=1'b1;
30342: pixelout<=1'b1;
30343: pixelout<=1'b1;
30344: pixelout<=1'b1;
30345: pixelout<=1'b1;
30346: pixelout<=1'b1;
30347: pixelout<=1'b1;
30348: pixelout<=1'b1;
30349: pixelout<=1'b1;
30350: pixelout<=1'b1;
30351: pixelout<=1'b1;
30352: pixelout<=1'b1;
30353: pixelout<=1'b1;
30354: pixelout<=1'b1;
30355: pixelout<=1'b1;
30356: pixelout<=1'b1;
30357: pixelout<=1'b1;
30358: pixelout<=1'b1;
30359: pixelout<=1'b1;
30360: pixelout<=1'b1;
30361: pixelout<=1'b1;
30362: pixelout<=1'b1;
30363: pixelout<=1'b1;
30364: pixelout<=1'b1;
30365: pixelout<=1'b1;
30366: pixelout<=1'b1;
30367: pixelout<=1'b1;
30368: pixelout<=1'b1;
30369: pixelout<=1'b1;
30370: pixelout<=1'b1;
30371: pixelout<=1'b1;
30372: pixelout<=1'b1;
30373: pixelout<=1'b1;
30374: pixelout<=1'b1;
30375: pixelout<=1'b1;
30376: pixelout<=1'b1;
30377: pixelout<=1'b1;
30378: pixelout<=1'b1;
30379: pixelout<=1'b1;
30380: pixelout<=1'b1;
30381: pixelout<=1'b1;
30382: pixelout<=1'b1;
30383: pixelout<=1'b1;
30384: pixelout<=1'b1;
30385: pixelout<=1'b1;
30386: pixelout<=1'b1;
30387: pixelout<=1'b1;
30388: pixelout<=1'b1;
30389: pixelout<=1'b1;
30390: pixelout<=1'b1;
30391: pixelout<=1'b1;
30392: pixelout<=1'b1;
30393: pixelout<=1'b1;
30394: pixelout<=1'b1;
30395: pixelout<=1'b1;
30396: pixelout<=1'b1;
30397: pixelout<=1'b1;
30398: pixelout<=1'b1;
30399: pixelout<=1'b1;
30400: pixelout<=1'b1;
30401: pixelout<=1'b1;
30402: pixelout<=1'b1;
30403: pixelout<=1'b1;
30404: pixelout<=1'b1;
30405: pixelout<=1'b1;
30406: pixelout<=1'b1;
30407: pixelout<=1'b1;
30408: pixelout<=1'b1;
30409: pixelout<=1'b1;
30410: pixelout<=1'b1;
30411: pixelout<=1'b1;
30412: pixelout<=1'b1;
30413: pixelout<=1'b1;
30414: pixelout<=1'b1;
30415: pixelout<=1'b1;
30416: pixelout<=1'b1;
30417: pixelout<=1'b1;
30418: pixelout<=1'b1;
30419: pixelout<=1'b1;
30420: pixelout<=1'b1;
30421: pixelout<=1'b1;
30422: pixelout<=1'b1;
30423: pixelout<=1'b1;
30424: pixelout<=1'b1;
30425: pixelout<=1'b1;
30426: pixelout<=1'b1;
30427: pixelout<=1'b1;
30428: pixelout<=1'b1;
30429: pixelout<=1'b1;
30430: pixelout<=1'b1;
30431: pixelout<=1'b1;
30432: pixelout<=1'b1;
30433: pixelout<=1'b1;
30434: pixelout<=1'b1;
30435: pixelout<=1'b1;
30436: pixelout<=1'b1;
30437: pixelout<=1'b1;
30438: pixelout<=1'b1;
30439: pixelout<=1'b1;
30440: pixelout<=1'b1;
30441: pixelout<=1'b1;
30442: pixelout<=1'b1;
30443: pixelout<=1'b1;
30444: pixelout<=1'b1;
30445: pixelout<=1'b1;
30446: pixelout<=1'b1;
30447: pixelout<=1'b1;
30448: pixelout<=1'b1;
30449: pixelout<=1'b1;
30450: pixelout<=1'b1;
30451: pixelout<=1'b1;
30452: pixelout<=1'b1;
30453: pixelout<=1'b1;
30454: pixelout<=1'b1;
30455: pixelout<=1'b1;
30456: pixelout<=1'b1;
30457: pixelout<=1'b1;
30458: pixelout<=1'b1;
30459: pixelout<=1'b1;
30460: pixelout<=1'b1;
30461: pixelout<=1'b1;
30462: pixelout<=1'b1;
30463: pixelout<=1'b1;
30464: pixelout<=1'b1;
30465: pixelout<=1'b1;
30466: pixelout<=1'b1;
30467: pixelout<=1'b1;
30468: pixelout<=1'b1;
30469: pixelout<=1'b1;
30470: pixelout<=1'b1;
30471: pixelout<=1'b1;
30472: pixelout<=1'b1;
30473: pixelout<=1'b1;
30474: pixelout<=1'b1;
30475: pixelout<=1'b1;
30476: pixelout<=1'b1;
30477: pixelout<=1'b1;
30478: pixelout<=1'b1;
30479: pixelout<=1'b1;
30480: pixelout<=1'b1;
30481: pixelout<=1'b1;
30482: pixelout<=1'b1;
30483: pixelout<=1'b1;
30484: pixelout<=1'b1;
30485: pixelout<=1'b1;
30486: pixelout<=1'b1;
30487: pixelout<=1'b1;
30488: pixelout<=1'b1;
30489: pixelout<=1'b1;
30490: pixelout<=1'b1;
30491: pixelout<=1'b1;
30492: pixelout<=1'b1;
30493: pixelout<=1'b1;
30494: pixelout<=1'b1;
30495: pixelout<=1'b1;
30496: pixelout<=1'b1;
30497: pixelout<=1'b1;
30498: pixelout<=1'b1;
30499: pixelout<=1'b1;
30500: pixelout<=1'b1;
30501: pixelout<=1'b1;
30502: pixelout<=1'b1;
30503: pixelout<=1'b1;
30504: pixelout<=1'b1;
30505: pixelout<=1'b1;
30506: pixelout<=1'b1;
30507: pixelout<=1'b1;
30508: pixelout<=1'b1;
30509: pixelout<=1'b1;
30510: pixelout<=1'b1;
30511: pixelout<=1'b1;
30512: pixelout<=1'b1;
30513: pixelout<=1'b1;
30514: pixelout<=1'b1;
30515: pixelout<=1'b1;
30516: pixelout<=1'b1;
30517: pixelout<=1'b1;
30518: pixelout<=1'b1;
30519: pixelout<=1'b1;
30520: pixelout<=1'b1;
30521: pixelout<=1'b1;
30522: pixelout<=1'b1;
30523: pixelout<=1'b1;
30524: pixelout<=1'b1;
30525: pixelout<=1'b1;
30526: pixelout<=1'b1;
30527: pixelout<=1'b1;
30528: pixelout<=1'b1;
30529: pixelout<=1'b1;
30530: pixelout<=1'b1;
30531: pixelout<=1'b1;
30532: pixelout<=1'b1;
30533: pixelout<=1'b1;
30534: pixelout<=1'b1;
30535: pixelout<=1'b1;
30536: pixelout<=1'b1;
30537: pixelout<=1'b1;
30538: pixelout<=1'b1;
30539: pixelout<=1'b1;
30540: pixelout<=1'b1;
30541: pixelout<=1'b1;
30542: pixelout<=1'b1;
30543: pixelout<=1'b1;
30544: pixelout<=1'b1;
30545: pixelout<=1'b1;
30546: pixelout<=1'b1;
30547: pixelout<=1'b1;
30548: pixelout<=1'b1;
30549: pixelout<=1'b1;
30550: pixelout<=1'b1;
30551: pixelout<=1'b1;
30552: pixelout<=1'b1;
30553: pixelout<=1'b1;
30554: pixelout<=1'b1;
30555: pixelout<=1'b1;
30556: pixelout<=1'b1;
30557: pixelout<=1'b1;
30558: pixelout<=1'b1;
30559: pixelout<=1'b1;
30560: pixelout<=1'b1;
30561: pixelout<=1'b1;
30562: pixelout<=1'b1;
30563: pixelout<=1'b1;
30564: pixelout<=1'b1;
30565: pixelout<=1'b1;
30566: pixelout<=1'b1;
30567: pixelout<=1'b1;
30568: pixelout<=1'b1;
30569: pixelout<=1'b1;
30570: pixelout<=1'b1;
30571: pixelout<=1'b1;
30572: pixelout<=1'b1;
30573: pixelout<=1'b1;
30574: pixelout<=1'b1;
30575: pixelout<=1'b1;
30576: pixelout<=1'b1;
30577: pixelout<=1'b1;
30578: pixelout<=1'b1;
30579: pixelout<=1'b1;
30580: pixelout<=1'b1;
30581: pixelout<=1'b1;
30582: pixelout<=1'b1;
30583: pixelout<=1'b1;
30584: pixelout<=1'b1;
30585: pixelout<=1'b1;
30586: pixelout<=1'b1;
30587: pixelout<=1'b1;
30588: pixelout<=1'b1;
30589: pixelout<=1'b1;
30590: pixelout<=1'b1;
30591: pixelout<=1'b1;
30592: pixelout<=1'b1;
30593: pixelout<=1'b1;
30594: pixelout<=1'b1;
30595: pixelout<=1'b1;
30596: pixelout<=1'b1;
30597: pixelout<=1'b1;
30598: pixelout<=1'b1;
30599: pixelout<=1'b1;
30600: pixelout<=1'b1;
30601: pixelout<=1'b1;
30602: pixelout<=1'b1;
30603: pixelout<=1'b1;
30604: pixelout<=1'b1;
30605: pixelout<=1'b1;
30606: pixelout<=1'b1;
30607: pixelout<=1'b1;
30608: pixelout<=1'b1;
30609: pixelout<=1'b1;
30610: pixelout<=1'b1;
30611: pixelout<=1'b1;
30612: pixelout<=1'b1;
30613: pixelout<=1'b1;
30614: pixelout<=1'b1;
30615: pixelout<=1'b1;
30616: pixelout<=1'b1;
30617: pixelout<=1'b1;
30618: pixelout<=1'b1;
30619: pixelout<=1'b1;
30620: pixelout<=1'b1;
30621: pixelout<=1'b1;
30622: pixelout<=1'b1;
30623: pixelout<=1'b1;
30624: pixelout<=1'b1;
30625: pixelout<=1'b1;
30626: pixelout<=1'b1;
30627: pixelout<=1'b1;
30628: pixelout<=1'b1;
30629: pixelout<=1'b1;
30630: pixelout<=1'b1;
30631: pixelout<=1'b1;
30632: pixelout<=1'b1;
30633: pixelout<=1'b1;
30634: pixelout<=1'b1;
30635: pixelout<=1'b1;
30636: pixelout<=1'b1;
30637: pixelout<=1'b1;
30638: pixelout<=1'b1;
30639: pixelout<=1'b1;
30640: pixelout<=1'b1;
30641: pixelout<=1'b1;
30642: pixelout<=1'b1;
30643: pixelout<=1'b1;
30644: pixelout<=1'b1;
30645: pixelout<=1'b1;
30646: pixelout<=1'b1;
30647: pixelout<=1'b1;
30648: pixelout<=1'b1;
30649: pixelout<=1'b1;
30650: pixelout<=1'b1;
30651: pixelout<=1'b1;
30652: pixelout<=1'b1;
30653: pixelout<=1'b1;
30654: pixelout<=1'b1;
30655: pixelout<=1'b1;
30656: pixelout<=1'b1;
30657: pixelout<=1'b1;
30658: pixelout<=1'b1;
30659: pixelout<=1'b1;
30660: pixelout<=1'b1;
30661: pixelout<=1'b1;
30662: pixelout<=1'b1;
30663: pixelout<=1'b1;
30664: pixelout<=1'b1;
30665: pixelout<=1'b1;
30666: pixelout<=1'b1;
30667: pixelout<=1'b1;
30668: pixelout<=1'b1;
30669: pixelout<=1'b1;
30670: pixelout<=1'b1;
30671: pixelout<=1'b1;
30672: pixelout<=1'b1;
30673: pixelout<=1'b1;
30674: pixelout<=1'b1;
30675: pixelout<=1'b1;
30676: pixelout<=1'b1;
30677: pixelout<=1'b1;
30678: pixelout<=1'b1;
30679: pixelout<=1'b1;
30680: pixelout<=1'b1;
30681: pixelout<=1'b1;
30682: pixelout<=1'b1;
30683: pixelout<=1'b1;
30684: pixelout<=1'b1;
30685: pixelout<=1'b1;
30686: pixelout<=1'b1;
30687: pixelout<=1'b1;
30688: pixelout<=1'b1;
30689: pixelout<=1'b1;
30690: pixelout<=1'b1;
30691: pixelout<=1'b1;
30692: pixelout<=1'b1;
30693: pixelout<=1'b1;
30694: pixelout<=1'b1;
30695: pixelout<=1'b1;
30696: pixelout<=1'b1;
30697: pixelout<=1'b1;
30698: pixelout<=1'b1;
30699: pixelout<=1'b1;
30700: pixelout<=1'b1;
30701: pixelout<=1'b1;
30702: pixelout<=1'b1;
30703: pixelout<=1'b1;
30704: pixelout<=1'b1;
30705: pixelout<=1'b1;
30706: pixelout<=1'b1;
30707: pixelout<=1'b1;
30708: pixelout<=1'b1;
30709: pixelout<=1'b1;
30710: pixelout<=1'b1;
30711: pixelout<=1'b1;
30712: pixelout<=1'b1;
30713: pixelout<=1'b1;
30714: pixelout<=1'b1;
30715: pixelout<=1'b1;
30716: pixelout<=1'b1;
30717: pixelout<=1'b1;
30718: pixelout<=1'b1;
30719: pixelout<=1'b1;
30720: pixelout<=1'b1;
30721: pixelout<=1'b1;
30722: pixelout<=1'b1;
30723: pixelout<=1'b1;
30724: pixelout<=1'b1;
30725: pixelout<=1'b1;
30726: pixelout<=1'b1;
30727: pixelout<=1'b1;
30728: pixelout<=1'b1;
30729: pixelout<=1'b1;
30730: pixelout<=1'b1;
30731: pixelout<=1'b1;
30732: pixelout<=1'b1;
30733: pixelout<=1'b1;
30734: pixelout<=1'b1;
30735: pixelout<=1'b1;
30736: pixelout<=1'b1;
30737: pixelout<=1'b1;
30738: pixelout<=1'b1;
30739: pixelout<=1'b1;
30740: pixelout<=1'b1;
30741: pixelout<=1'b1;
30742: pixelout<=1'b1;
30743: pixelout<=1'b1;
30744: pixelout<=1'b1;
30745: pixelout<=1'b1;
30746: pixelout<=1'b1;
30747: pixelout<=1'b1;
30748: pixelout<=1'b1;
30749: pixelout<=1'b1;
30750: pixelout<=1'b1;
30751: pixelout<=1'b1;
30752: pixelout<=1'b1;
30753: pixelout<=1'b1;
30754: pixelout<=1'b1;
30755: pixelout<=1'b1;
30756: pixelout<=1'b1;
30757: pixelout<=1'b1;
30758: pixelout<=1'b1;
30759: pixelout<=1'b1;
30760: pixelout<=1'b1;
30761: pixelout<=1'b1;
30762: pixelout<=1'b1;
30763: pixelout<=1'b1;
30764: pixelout<=1'b1;
30765: pixelout<=1'b1;
30766: pixelout<=1'b1;
30767: pixelout<=1'b1;
30768: pixelout<=1'b1;
30769: pixelout<=1'b1;
30770: pixelout<=1'b1;
30771: pixelout<=1'b1;
30772: pixelout<=1'b1;
30773: pixelout<=1'b1;
30774: pixelout<=1'b1;
30775: pixelout<=1'b1;
30776: pixelout<=1'b1;
30777: pixelout<=1'b1;
30778: pixelout<=1'b1;
30779: pixelout<=1'b1;
30780: pixelout<=1'b1;
30781: pixelout<=1'b1;
30782: pixelout<=1'b1;
30783: pixelout<=1'b1;
30784: pixelout<=1'b1;
30785: pixelout<=1'b1;
30786: pixelout<=1'b1;
30787: pixelout<=1'b1;
30788: pixelout<=1'b1;
30789: pixelout<=1'b1;
30790: pixelout<=1'b1;
30791: pixelout<=1'b1;
30792: pixelout<=1'b1;
30793: pixelout<=1'b1;
30794: pixelout<=1'b1;
30795: pixelout<=1'b1;
30796: pixelout<=1'b1;
30797: pixelout<=1'b1;
30798: pixelout<=1'b1;
30799: pixelout<=1'b1;
30800: pixelout<=1'b1;
30801: pixelout<=1'b1;
30802: pixelout<=1'b1;
30803: pixelout<=1'b1;
30804: pixelout<=1'b1;
30805: pixelout<=1'b1;
30806: pixelout<=1'b1;
30807: pixelout<=1'b1;
30808: pixelout<=1'b1;
30809: pixelout<=1'b1;
30810: pixelout<=1'b1;
30811: pixelout<=1'b1;
30812: pixelout<=1'b1;
30813: pixelout<=1'b1;
30814: pixelout<=1'b1;
30815: pixelout<=1'b1;
30816: pixelout<=1'b1;
30817: pixelout<=1'b1;
30818: pixelout<=1'b1;
30819: pixelout<=1'b1;
30820: pixelout<=1'b1;
30821: pixelout<=1'b1;
30822: pixelout<=1'b1;
30823: pixelout<=1'b1;
30824: pixelout<=1'b1;
30825: pixelout<=1'b1;
30826: pixelout<=1'b1;
30827: pixelout<=1'b1;
30828: pixelout<=1'b1;
30829: pixelout<=1'b1;
30830: pixelout<=1'b1;
30831: pixelout<=1'b1;
30832: pixelout<=1'b1;
30833: pixelout<=1'b1;
30834: pixelout<=1'b1;
30835: pixelout<=1'b1;
30836: pixelout<=1'b1;
30837: pixelout<=1'b1;
30838: pixelout<=1'b1;
30839: pixelout<=1'b1;
30840: pixelout<=1'b1;
30841: pixelout<=1'b1;
30842: pixelout<=1'b1;
30843: pixelout<=1'b1;
30844: pixelout<=1'b1;
30845: pixelout<=1'b1;
30846: pixelout<=1'b1;
30847: pixelout<=1'b1;
30848: pixelout<=1'b1;
30849: pixelout<=1'b1;
30850: pixelout<=1'b1;
30851: pixelout<=1'b1;
30852: pixelout<=1'b1;
30853: pixelout<=1'b1;
30854: pixelout<=1'b1;
30855: pixelout<=1'b1;
30856: pixelout<=1'b1;
30857: pixelout<=1'b1;
30858: pixelout<=1'b1;
30859: pixelout<=1'b1;
30860: pixelout<=1'b1;
30861: pixelout<=1'b1;
30862: pixelout<=1'b1;
30863: pixelout<=1'b1;
30864: pixelout<=1'b1;
30865: pixelout<=1'b1;
30866: pixelout<=1'b1;
30867: pixelout<=1'b1;
30868: pixelout<=1'b1;
30869: pixelout<=1'b1;
30870: pixelout<=1'b1;
30871: pixelout<=1'b1;
30872: pixelout<=1'b1;
30873: pixelout<=1'b1;
30874: pixelout<=1'b1;
30875: pixelout<=1'b1;
30876: pixelout<=1'b1;
30877: pixelout<=1'b1;
30878: pixelout<=1'b1;
30879: pixelout<=1'b1;
30880: pixelout<=1'b1;
30881: pixelout<=1'b1;
30882: pixelout<=1'b1;
30883: pixelout<=1'b1;
30884: pixelout<=1'b1;
30885: pixelout<=1'b1;
30886: pixelout<=1'b1;
30887: pixelout<=1'b1;
30888: pixelout<=1'b1;
30889: pixelout<=1'b1;
30890: pixelout<=1'b1;
30891: pixelout<=1'b1;
30892: pixelout<=1'b1;
30893: pixelout<=1'b1;
30894: pixelout<=1'b1;
30895: pixelout<=1'b1;
30896: pixelout<=1'b1;
30897: pixelout<=1'b1;
30898: pixelout<=1'b1;
30899: pixelout<=1'b1;
30900: pixelout<=1'b1;
30901: pixelout<=1'b1;
30902: pixelout<=1'b1;
30903: pixelout<=1'b1;
30904: pixelout<=1'b1;
30905: pixelout<=1'b1;
30906: pixelout<=1'b1;
30907: pixelout<=1'b1;
30908: pixelout<=1'b1;
30909: pixelout<=1'b1;
30910: pixelout<=1'b1;
30911: pixelout<=1'b1;
30912: pixelout<=1'b1;
30913: pixelout<=1'b1;
30914: pixelout<=1'b1;
30915: pixelout<=1'b1;
30916: pixelout<=1'b1;
30917: pixelout<=1'b1;
30918: pixelout<=1'b1;
30919: pixelout<=1'b1;
30920: pixelout<=1'b1;
30921: pixelout<=1'b1;
30922: pixelout<=1'b1;
30923: pixelout<=1'b1;
30924: pixelout<=1'b1;
30925: pixelout<=1'b1;
30926: pixelout<=1'b1;
30927: pixelout<=1'b1;
30928: pixelout<=1'b1;
30929: pixelout<=1'b1;
30930: pixelout<=1'b1;
30931: pixelout<=1'b1;
30932: pixelout<=1'b1;
30933: pixelout<=1'b1;
30934: pixelout<=1'b1;
30935: pixelout<=1'b1;
30936: pixelout<=1'b1;
30937: pixelout<=1'b1;
30938: pixelout<=1'b1;
30939: pixelout<=1'b1;
30940: pixelout<=1'b1;
30941: pixelout<=1'b1;
30942: pixelout<=1'b1;
30943: pixelout<=1'b1;
30944: pixelout<=1'b1;
30945: pixelout<=1'b1;
30946: pixelout<=1'b1;
30947: pixelout<=1'b1;
30948: pixelout<=1'b1;
30949: pixelout<=1'b1;
30950: pixelout<=1'b1;
30951: pixelout<=1'b1;
30952: pixelout<=1'b1;
30953: pixelout<=1'b1;
30954: pixelout<=1'b1;
30955: pixelout<=1'b1;
30956: pixelout<=1'b1;
30957: pixelout<=1'b1;
30958: pixelout<=1'b1;
30959: pixelout<=1'b1;
30960: pixelout<=1'b1;
30961: pixelout<=1'b1;
30962: pixelout<=1'b1;
30963: pixelout<=1'b1;
30964: pixelout<=1'b1;
30965: pixelout<=1'b1;
30966: pixelout<=1'b1;
30967: pixelout<=1'b1;
30968: pixelout<=1'b1;
30969: pixelout<=1'b1;
30970: pixelout<=1'b1;
30971: pixelout<=1'b1;
30972: pixelout<=1'b1;
30973: pixelout<=1'b1;
30974: pixelout<=1'b1;
30975: pixelout<=1'b1;
30976: pixelout<=1'b1;
30977: pixelout<=1'b1;
30978: pixelout<=1'b1;
30979: pixelout<=1'b1;
30980: pixelout<=1'b1;
30981: pixelout<=1'b1;
30982: pixelout<=1'b1;
30983: pixelout<=1'b1;
30984: pixelout<=1'b1;
30985: pixelout<=1'b1;
30986: pixelout<=1'b1;
30987: pixelout<=1'b1;
30988: pixelout<=1'b1;
30989: pixelout<=1'b1;
30990: pixelout<=1'b1;
30991: pixelout<=1'b1;
30992: pixelout<=1'b1;
30993: pixelout<=1'b1;
30994: pixelout<=1'b1;
30995: pixelout<=1'b1;
30996: pixelout<=1'b1;
30997: pixelout<=1'b1;
30998: pixelout<=1'b1;
30999: pixelout<=1'b1;
31000: pixelout<=1'b1;
31001: pixelout<=1'b1;
31002: pixelout<=1'b1;
31003: pixelout<=1'b1;
31004: pixelout<=1'b1;
31005: pixelout<=1'b1;
31006: pixelout<=1'b1;
31007: pixelout<=1'b1;
31008: pixelout<=1'b1;
31009: pixelout<=1'b1;
31010: pixelout<=1'b1;
31011: pixelout<=1'b1;
31012: pixelout<=1'b1;
31013: pixelout<=1'b1;
31014: pixelout<=1'b1;
31015: pixelout<=1'b1;
31016: pixelout<=1'b1;
31017: pixelout<=1'b1;
31018: pixelout<=1'b1;
31019: pixelout<=1'b1;
31020: pixelout<=1'b1;
31021: pixelout<=1'b1;
31022: pixelout<=1'b1;
31023: pixelout<=1'b1;
31024: pixelout<=1'b1;
31025: pixelout<=1'b1;
31026: pixelout<=1'b1;
31027: pixelout<=1'b1;
31028: pixelout<=1'b1;
31029: pixelout<=1'b1;
31030: pixelout<=1'b1;
31031: pixelout<=1'b1;
31032: pixelout<=1'b1;
31033: pixelout<=1'b1;
31034: pixelout<=1'b1;
31035: pixelout<=1'b1;
31036: pixelout<=1'b1;
31037: pixelout<=1'b1;
31038: pixelout<=1'b1;
31039: pixelout<=1'b1;
31040: pixelout<=1'b1;
31041: pixelout<=1'b1;
31042: pixelout<=1'b1;
31043: pixelout<=1'b1;
31044: pixelout<=1'b1;
31045: pixelout<=1'b1;
31046: pixelout<=1'b1;
31047: pixelout<=1'b1;
31048: pixelout<=1'b1;
31049: pixelout<=1'b1;
31050: pixelout<=1'b1;
31051: pixelout<=1'b1;
31052: pixelout<=1'b1;
31053: pixelout<=1'b1;
31054: pixelout<=1'b1;
31055: pixelout<=1'b1;
31056: pixelout<=1'b1;
31057: pixelout<=1'b1;
31058: pixelout<=1'b1;
31059: pixelout<=1'b1;
31060: pixelout<=1'b1;
31061: pixelout<=1'b1;
31062: pixelout<=1'b1;
31063: pixelout<=1'b1;
31064: pixelout<=1'b1;
31065: pixelout<=1'b1;
31066: pixelout<=1'b1;
31067: pixelout<=1'b1;
31068: pixelout<=1'b1;
31069: pixelout<=1'b1;
31070: pixelout<=1'b1;
31071: pixelout<=1'b1;
31072: pixelout<=1'b1;
31073: pixelout<=1'b1;
31074: pixelout<=1'b1;
31075: pixelout<=1'b1;
31076: pixelout<=1'b1;
31077: pixelout<=1'b1;
31078: pixelout<=1'b1;
31079: pixelout<=1'b1;
31080: pixelout<=1'b1;
31081: pixelout<=1'b1;
31082: pixelout<=1'b1;
31083: pixelout<=1'b1;
31084: pixelout<=1'b1;
31085: pixelout<=1'b1;
31086: pixelout<=1'b1;
31087: pixelout<=1'b1;
31088: pixelout<=1'b1;
31089: pixelout<=1'b1;
31090: pixelout<=1'b1;
31091: pixelout<=1'b1;
31092: pixelout<=1'b1;
31093: pixelout<=1'b1;
31094: pixelout<=1'b1;
31095: pixelout<=1'b1;
31096: pixelout<=1'b1;
31097: pixelout<=1'b1;
31098: pixelout<=1'b1;
31099: pixelout<=1'b1;
31100: pixelout<=1'b1;
31101: pixelout<=1'b1;
31102: pixelout<=1'b1;
31103: pixelout<=1'b1;
31104: pixelout<=1'b1;
31105: pixelout<=1'b1;
31106: pixelout<=1'b1;
31107: pixelout<=1'b1;
31108: pixelout<=1'b1;
31109: pixelout<=1'b1;
31110: pixelout<=1'b1;
31111: pixelout<=1'b1;
31112: pixelout<=1'b1;
31113: pixelout<=1'b1;
31114: pixelout<=1'b1;
31115: pixelout<=1'b1;
31116: pixelout<=1'b1;
31117: pixelout<=1'b1;
31118: pixelout<=1'b1;
31119: pixelout<=1'b1;
31120: pixelout<=1'b1;
31121: pixelout<=1'b1;
31122: pixelout<=1'b1;
31123: pixelout<=1'b1;
31124: pixelout<=1'b1;
31125: pixelout<=1'b1;
31126: pixelout<=1'b1;
31127: pixelout<=1'b1;
31128: pixelout<=1'b1;
31129: pixelout<=1'b1;
31130: pixelout<=1'b1;
31131: pixelout<=1'b1;
31132: pixelout<=1'b1;
31133: pixelout<=1'b1;
31134: pixelout<=1'b1;
31135: pixelout<=1'b1;
31136: pixelout<=1'b1;
31137: pixelout<=1'b1;
31138: pixelout<=1'b1;
31139: pixelout<=1'b1;
31140: pixelout<=1'b1;
31141: pixelout<=1'b1;
31142: pixelout<=1'b1;
31143: pixelout<=1'b1;
31144: pixelout<=1'b1;
31145: pixelout<=1'b1;
31146: pixelout<=1'b1;
31147: pixelout<=1'b1;
31148: pixelout<=1'b1;
31149: pixelout<=1'b1;
31150: pixelout<=1'b1;
31151: pixelout<=1'b1;
31152: pixelout<=1'b1;
31153: pixelout<=1'b1;
31154: pixelout<=1'b1;
31155: pixelout<=1'b1;
31156: pixelout<=1'b1;
31157: pixelout<=1'b1;
31158: pixelout<=1'b1;
31159: pixelout<=1'b1;
31160: pixelout<=1'b1;
31161: pixelout<=1'b1;
31162: pixelout<=1'b1;
31163: pixelout<=1'b1;
31164: pixelout<=1'b1;
31165: pixelout<=1'b1;
31166: pixelout<=1'b1;
31167: pixelout<=1'b1;
31168: pixelout<=1'b1;
31169: pixelout<=1'b1;
31170: pixelout<=1'b1;
31171: pixelout<=1'b1;
31172: pixelout<=1'b1;
31173: pixelout<=1'b1;
31174: pixelout<=1'b1;
31175: pixelout<=1'b1;
31176: pixelout<=1'b1;
31177: pixelout<=1'b1;
31178: pixelout<=1'b1;
31179: pixelout<=1'b1;
31180: pixelout<=1'b1;
31181: pixelout<=1'b1;
31182: pixelout<=1'b1;
31183: pixelout<=1'b1;
31184: pixelout<=1'b1;
31185: pixelout<=1'b1;
31186: pixelout<=1'b1;
31187: pixelout<=1'b1;
31188: pixelout<=1'b1;
31189: pixelout<=1'b1;
31190: pixelout<=1'b1;
31191: pixelout<=1'b1;
31192: pixelout<=1'b1;
31193: pixelout<=1'b1;
31194: pixelout<=1'b1;
31195: pixelout<=1'b1;
31196: pixelout<=1'b1;
31197: pixelout<=1'b1;
31198: pixelout<=1'b1;
31199: pixelout<=1'b1;
31200: pixelout<=1'b1;
31201: pixelout<=1'b1;
31202: pixelout<=1'b1;
31203: pixelout<=1'b1;
31204: pixelout<=1'b1;
31205: pixelout<=1'b1;
31206: pixelout<=1'b1;
31207: pixelout<=1'b1;
31208: pixelout<=1'b1;
31209: pixelout<=1'b1;
31210: pixelout<=1'b1;
31211: pixelout<=1'b1;
31212: pixelout<=1'b1;
31213: pixelout<=1'b1;
31214: pixelout<=1'b1;
31215: pixelout<=1'b1;
31216: pixelout<=1'b1;
31217: pixelout<=1'b1;
31218: pixelout<=1'b1;
31219: pixelout<=1'b1;
31220: pixelout<=1'b1;
31221: pixelout<=1'b1;
31222: pixelout<=1'b1;
31223: pixelout<=1'b1;
31224: pixelout<=1'b1;
31225: pixelout<=1'b1;
31226: pixelout<=1'b1;
31227: pixelout<=1'b1;
31228: pixelout<=1'b1;
31229: pixelout<=1'b1;
31230: pixelout<=1'b1;
31231: pixelout<=1'b1;
31232: pixelout<=1'b1;
31233: pixelout<=1'b1;
31234: pixelout<=1'b1;
31235: pixelout<=1'b1;
31236: pixelout<=1'b1;
31237: pixelout<=1'b1;
31238: pixelout<=1'b1;
31239: pixelout<=1'b1;
31240: pixelout<=1'b1;
31241: pixelout<=1'b1;
31242: pixelout<=1'b1;
31243: pixelout<=1'b1;
31244: pixelout<=1'b1;
31245: pixelout<=1'b1;
31246: pixelout<=1'b1;
31247: pixelout<=1'b1;
31248: pixelout<=1'b1;
31249: pixelout<=1'b1;
31250: pixelout<=1'b1;
31251: pixelout<=1'b1;
31252: pixelout<=1'b1;
31253: pixelout<=1'b1;
31254: pixelout<=1'b1;
31255: pixelout<=1'b1;
31256: pixelout<=1'b1;
31257: pixelout<=1'b1;
31258: pixelout<=1'b1;
31259: pixelout<=1'b1;
31260: pixelout<=1'b1;
31261: pixelout<=1'b1;
31262: pixelout<=1'b1;
31263: pixelout<=1'b1;
31264: pixelout<=1'b1;
31265: pixelout<=1'b1;
31266: pixelout<=1'b1;
31267: pixelout<=1'b1;
31268: pixelout<=1'b1;
31269: pixelout<=1'b1;
31270: pixelout<=1'b1;
31271: pixelout<=1'b1;
31272: pixelout<=1'b1;
31273: pixelout<=1'b1;
31274: pixelout<=1'b1;
31275: pixelout<=1'b1;
31276: pixelout<=1'b1;
31277: pixelout<=1'b1;
31278: pixelout<=1'b1;
31279: pixelout<=1'b1;
31280: pixelout<=1'b1;
31281: pixelout<=1'b1;
31282: pixelout<=1'b1;
31283: pixelout<=1'b1;
31284: pixelout<=1'b1;
31285: pixelout<=1'b1;
31286: pixelout<=1'b1;
31287: pixelout<=1'b1;
31288: pixelout<=1'b1;
31289: pixelout<=1'b1;
31290: pixelout<=1'b1;
31291: pixelout<=1'b1;
31292: pixelout<=1'b1;
31293: pixelout<=1'b1;
31294: pixelout<=1'b1;
31295: pixelout<=1'b1;
31296: pixelout<=1'b1;
31297: pixelout<=1'b1;
31298: pixelout<=1'b1;
31299: pixelout<=1'b1;
31300: pixelout<=1'b1;
31301: pixelout<=1'b1;
31302: pixelout<=1'b1;
31303: pixelout<=1'b1;
31304: pixelout<=1'b1;
31305: pixelout<=1'b1;
31306: pixelout<=1'b1;
31307: pixelout<=1'b1;
31308: pixelout<=1'b1;
31309: pixelout<=1'b1;
31310: pixelout<=1'b1;
31311: pixelout<=1'b1;
31312: pixelout<=1'b1;
31313: pixelout<=1'b1;
31314: pixelout<=1'b1;
31315: pixelout<=1'b1;
31316: pixelout<=1'b1;
31317: pixelout<=1'b1;
31318: pixelout<=1'b1;
31319: pixelout<=1'b1;
31320: pixelout<=1'b1;
31321: pixelout<=1'b1;
31322: pixelout<=1'b1;
31323: pixelout<=1'b1;
31324: pixelout<=1'b1;
31325: pixelout<=1'b1;
31326: pixelout<=1'b1;
31327: pixelout<=1'b1;
31328: pixelout<=1'b1;
31329: pixelout<=1'b1;
31330: pixelout<=1'b0;
31331: pixelout<=1'b0;
31332: pixelout<=1'b0;
31333: pixelout<=1'b1;
31334: pixelout<=1'b1;
31335: pixelout<=1'b1;
31336: pixelout<=1'b1;
31337: pixelout<=1'b1;
31338: pixelout<=1'b1;
31339: pixelout<=1'b1;
31340: pixelout<=1'b1;
31341: pixelout<=1'b1;
31342: pixelout<=1'b1;
31343: pixelout<=1'b1;
31344: pixelout<=1'b1;
31345: pixelout<=1'b1;
31346: pixelout<=1'b1;
31347: pixelout<=1'b1;
31348: pixelout<=1'b1;
31349: pixelout<=1'b1;
31350: pixelout<=1'b1;
31351: pixelout<=1'b1;
31352: pixelout<=1'b1;
31353: pixelout<=1'b1;
31354: pixelout<=1'b1;
31355: pixelout<=1'b1;
31356: pixelout<=1'b1;
31357: pixelout<=1'b1;
31358: pixelout<=1'b1;
31359: pixelout<=1'b1;
31360: pixelout<=1'b1;
31361: pixelout<=1'b1;
31362: pixelout<=1'b1;
31363: pixelout<=1'b1;
31364: pixelout<=1'b1;
31365: pixelout<=1'b1;
31366: pixelout<=1'b1;
31367: pixelout<=1'b1;
31368: pixelout<=1'b1;
31369: pixelout<=1'b1;
31370: pixelout<=1'b1;
31371: pixelout<=1'b0;
31372: pixelout<=1'b1;
31373: pixelout<=1'b1;
31374: pixelout<=1'b1;
31375: pixelout<=1'b0;
31376: pixelout<=1'b0;
31377: pixelout<=1'b0;
31378: pixelout<=1'b0;
31379: pixelout<=1'b0;
31380: pixelout<=1'b1;
31381: pixelout<=1'b1;
31382: pixelout<=1'b1;
31383: pixelout<=1'b1;
31384: pixelout<=1'b1;
31385: pixelout<=1'b1;
31386: pixelout<=1'b1;
31387: pixelout<=1'b1;
31388: pixelout<=1'b1;
31389: pixelout<=1'b1;
31390: pixelout<=1'b0;
31391: pixelout<=1'b1;
31392: pixelout<=1'b1;
31393: pixelout<=1'b1;
31394: pixelout<=1'b1;
31395: pixelout<=1'b1;
31396: pixelout<=1'b1;
31397: pixelout<=1'b1;
31398: pixelout<=1'b1;
31399: pixelout<=1'b1;
31400: pixelout<=1'b1;
31401: pixelout<=1'b1;
31402: pixelout<=1'b1;
31403: pixelout<=1'b1;
31404: pixelout<=1'b1;
31405: pixelout<=1'b1;
31406: pixelout<=1'b1;
31407: pixelout<=1'b1;
31408: pixelout<=1'b1;
31409: pixelout<=1'b1;
31410: pixelout<=1'b1;
31411: pixelout<=1'b1;
31412: pixelout<=1'b1;
31413: pixelout<=1'b1;
31414: pixelout<=1'b1;
31415: pixelout<=1'b1;
31416: pixelout<=1'b1;
31417: pixelout<=1'b1;
31418: pixelout<=1'b1;
31419: pixelout<=1'b1;
31420: pixelout<=1'b1;
31421: pixelout<=1'b1;
31422: pixelout<=1'b1;
31423: pixelout<=1'b1;
31424: pixelout<=1'b1;
31425: pixelout<=1'b1;
31426: pixelout<=1'b1;
31427: pixelout<=1'b1;
31428: pixelout<=1'b1;
31429: pixelout<=1'b1;
31430: pixelout<=1'b1;
31431: pixelout<=1'b1;
31432: pixelout<=1'b1;
31433: pixelout<=1'b1;
31434: pixelout<=1'b1;
31435: pixelout<=1'b1;
31436: pixelout<=1'b1;
31437: pixelout<=1'b1;
31438: pixelout<=1'b1;
31439: pixelout<=1'b1;
31440: pixelout<=1'b1;
31441: pixelout<=1'b1;
31442: pixelout<=1'b1;
31443: pixelout<=1'b1;
31444: pixelout<=1'b1;
31445: pixelout<=1'b1;
31446: pixelout<=1'b1;
31447: pixelout<=1'b1;
31448: pixelout<=1'b1;
31449: pixelout<=1'b1;
31450: pixelout<=1'b1;
31451: pixelout<=1'b1;
31452: pixelout<=1'b1;
31453: pixelout<=1'b1;
31454: pixelout<=1'b1;
31455: pixelout<=1'b1;
31456: pixelout<=1'b1;
31457: pixelout<=1'b1;
31458: pixelout<=1'b1;
31459: pixelout<=1'b1;
31460: pixelout<=1'b1;
31461: pixelout<=1'b1;
31462: pixelout<=1'b1;
31463: pixelout<=1'b1;
31464: pixelout<=1'b1;
31465: pixelout<=1'b1;
31466: pixelout<=1'b1;
31467: pixelout<=1'b1;
31468: pixelout<=1'b1;
31469: pixelout<=1'b1;
31470: pixelout<=1'b1;
31471: pixelout<=1'b1;
31472: pixelout<=1'b1;
31473: pixelout<=1'b1;
31474: pixelout<=1'b1;
31475: pixelout<=1'b1;
31476: pixelout<=1'b1;
31477: pixelout<=1'b1;
31478: pixelout<=1'b1;
31479: pixelout<=1'b1;
31480: pixelout<=1'b1;
31481: pixelout<=1'b1;
31482: pixelout<=1'b1;
31483: pixelout<=1'b1;
31484: pixelout<=1'b1;
31485: pixelout<=1'b1;
31486: pixelout<=1'b1;
31487: pixelout<=1'b1;
31488: pixelout<=1'b1;
31489: pixelout<=1'b1;
31490: pixelout<=1'b1;
31491: pixelout<=1'b1;
31492: pixelout<=1'b1;
31493: pixelout<=1'b1;
31494: pixelout<=1'b1;
31495: pixelout<=1'b1;
31496: pixelout<=1'b1;
31497: pixelout<=1'b1;
31498: pixelout<=1'b1;
31499: pixelout<=1'b1;
31500: pixelout<=1'b1;
31501: pixelout<=1'b1;
31502: pixelout<=1'b1;
31503: pixelout<=1'b1;
31504: pixelout<=1'b1;
31505: pixelout<=1'b1;
31506: pixelout<=1'b1;
31507: pixelout<=1'b1;
31508: pixelout<=1'b1;
31509: pixelout<=1'b1;
31510: pixelout<=1'b1;
31511: pixelout<=1'b1;
31512: pixelout<=1'b1;
31513: pixelout<=1'b1;
31514: pixelout<=1'b1;
31515: pixelout<=1'b0;
31516: pixelout<=1'b1;
31517: pixelout<=1'b1;
31518: pixelout<=1'b1;
31519: pixelout<=1'b1;
31520: pixelout<=1'b1;
31521: pixelout<=1'b1;
31522: pixelout<=1'b1;
31523: pixelout<=1'b1;
31524: pixelout<=1'b1;
31525: pixelout<=1'b1;
31526: pixelout<=1'b1;
31527: pixelout<=1'b1;
31528: pixelout<=1'b1;
31529: pixelout<=1'b1;
31530: pixelout<=1'b1;
31531: pixelout<=1'b1;
31532: pixelout<=1'b1;
31533: pixelout<=1'b1;
31534: pixelout<=1'b1;
31535: pixelout<=1'b1;
31536: pixelout<=1'b1;
31537: pixelout<=1'b1;
31538: pixelout<=1'b1;
31539: pixelout<=1'b1;
31540: pixelout<=1'b1;
31541: pixelout<=1'b1;
31542: pixelout<=1'b1;
31543: pixelout<=1'b1;
31544: pixelout<=1'b1;
31545: pixelout<=1'b1;
31546: pixelout<=1'b1;
31547: pixelout<=1'b1;
31548: pixelout<=1'b1;
31549: pixelout<=1'b1;
31550: pixelout<=1'b1;
31551: pixelout<=1'b1;
31552: pixelout<=1'b1;
31553: pixelout<=1'b1;
31554: pixelout<=1'b1;
31555: pixelout<=1'b1;
31556: pixelout<=1'b1;
31557: pixelout<=1'b1;
31558: pixelout<=1'b1;
31559: pixelout<=1'b1;
31560: pixelout<=1'b1;
31561: pixelout<=1'b1;
31562: pixelout<=1'b1;
31563: pixelout<=1'b1;
31564: pixelout<=1'b1;
31565: pixelout<=1'b1;
31566: pixelout<=1'b1;
31567: pixelout<=1'b1;
31568: pixelout<=1'b1;
31569: pixelout<=1'b0;
31570: pixelout<=1'b1;
31571: pixelout<=1'b1;
31572: pixelout<=1'b1;
31573: pixelout<=1'b0;
31574: pixelout<=1'b1;
31575: pixelout<=1'b1;
31576: pixelout<=1'b1;
31577: pixelout<=1'b1;
31578: pixelout<=1'b1;
31579: pixelout<=1'b1;
31580: pixelout<=1'b1;
31581: pixelout<=1'b1;
31582: pixelout<=1'b1;
31583: pixelout<=1'b1;
31584: pixelout<=1'b1;
31585: pixelout<=1'b1;
31586: pixelout<=1'b1;
31587: pixelout<=1'b1;
31588: pixelout<=1'b1;
31589: pixelout<=1'b1;
31590: pixelout<=1'b1;
31591: pixelout<=1'b1;
31592: pixelout<=1'b1;
31593: pixelout<=1'b1;
31594: pixelout<=1'b1;
31595: pixelout<=1'b1;
31596: pixelout<=1'b1;
31597: pixelout<=1'b1;
31598: pixelout<=1'b1;
31599: pixelout<=1'b1;
31600: pixelout<=1'b1;
31601: pixelout<=1'b1;
31602: pixelout<=1'b1;
31603: pixelout<=1'b1;
31604: pixelout<=1'b1;
31605: pixelout<=1'b1;
31606: pixelout<=1'b1;
31607: pixelout<=1'b1;
31608: pixelout<=1'b1;
31609: pixelout<=1'b1;
31610: pixelout<=1'b1;
31611: pixelout<=1'b0;
31612: pixelout<=1'b1;
31613: pixelout<=1'b1;
31614: pixelout<=1'b1;
31615: pixelout<=1'b0;
31616: pixelout<=1'b1;
31617: pixelout<=1'b1;
31618: pixelout<=1'b1;
31619: pixelout<=1'b1;
31620: pixelout<=1'b1;
31621: pixelout<=1'b1;
31622: pixelout<=1'b1;
31623: pixelout<=1'b1;
31624: pixelout<=1'b1;
31625: pixelout<=1'b1;
31626: pixelout<=1'b1;
31627: pixelout<=1'b1;
31628: pixelout<=1'b1;
31629: pixelout<=1'b1;
31630: pixelout<=1'b0;
31631: pixelout<=1'b1;
31632: pixelout<=1'b1;
31633: pixelout<=1'b1;
31634: pixelout<=1'b1;
31635: pixelout<=1'b1;
31636: pixelout<=1'b1;
31637: pixelout<=1'b1;
31638: pixelout<=1'b1;
31639: pixelout<=1'b1;
31640: pixelout<=1'b1;
31641: pixelout<=1'b1;
31642: pixelout<=1'b1;
31643: pixelout<=1'b1;
31644: pixelout<=1'b1;
31645: pixelout<=1'b1;
31646: pixelout<=1'b1;
31647: pixelout<=1'b1;
31648: pixelout<=1'b1;
31649: pixelout<=1'b1;
31650: pixelout<=1'b1;
31651: pixelout<=1'b1;
31652: pixelout<=1'b1;
31653: pixelout<=1'b1;
31654: pixelout<=1'b1;
31655: pixelout<=1'b1;
31656: pixelout<=1'b1;
31657: pixelout<=1'b1;
31658: pixelout<=1'b1;
31659: pixelout<=1'b1;
31660: pixelout<=1'b1;
31661: pixelout<=1'b1;
31662: pixelout<=1'b1;
31663: pixelout<=1'b1;
31664: pixelout<=1'b1;
31665: pixelout<=1'b1;
31666: pixelout<=1'b1;
31667: pixelout<=1'b1;
31668: pixelout<=1'b1;
31669: pixelout<=1'b1;
31670: pixelout<=1'b1;
31671: pixelout<=1'b1;
31672: pixelout<=1'b1;
31673: pixelout<=1'b1;
31674: pixelout<=1'b1;
31675: pixelout<=1'b1;
31676: pixelout<=1'b1;
31677: pixelout<=1'b1;
31678: pixelout<=1'b1;
31679: pixelout<=1'b1;
31680: pixelout<=1'b1;
31681: pixelout<=1'b1;
31682: pixelout<=1'b1;
31683: pixelout<=1'b1;
31684: pixelout<=1'b1;
31685: pixelout<=1'b1;
31686: pixelout<=1'b1;
31687: pixelout<=1'b1;
31688: pixelout<=1'b1;
31689: pixelout<=1'b1;
31690: pixelout<=1'b1;
31691: pixelout<=1'b1;
31692: pixelout<=1'b1;
31693: pixelout<=1'b1;
31694: pixelout<=1'b1;
31695: pixelout<=1'b1;
31696: pixelout<=1'b1;
31697: pixelout<=1'b1;
31698: pixelout<=1'b1;
31699: pixelout<=1'b1;
31700: pixelout<=1'b1;
31701: pixelout<=1'b1;
31702: pixelout<=1'b1;
31703: pixelout<=1'b1;
31704: pixelout<=1'b1;
31705: pixelout<=1'b1;
31706: pixelout<=1'b1;
31707: pixelout<=1'b1;
31708: pixelout<=1'b1;
31709: pixelout<=1'b1;
31710: pixelout<=1'b1;
31711: pixelout<=1'b1;
31712: pixelout<=1'b1;
31713: pixelout<=1'b1;
31714: pixelout<=1'b1;
31715: pixelout<=1'b1;
31716: pixelout<=1'b1;
31717: pixelout<=1'b1;
31718: pixelout<=1'b1;
31719: pixelout<=1'b1;
31720: pixelout<=1'b1;
31721: pixelout<=1'b1;
31722: pixelout<=1'b1;
31723: pixelout<=1'b1;
31724: pixelout<=1'b1;
31725: pixelout<=1'b1;
31726: pixelout<=1'b1;
31727: pixelout<=1'b1;
31728: pixelout<=1'b1;
31729: pixelout<=1'b1;
31730: pixelout<=1'b1;
31731: pixelout<=1'b1;
31732: pixelout<=1'b1;
31733: pixelout<=1'b1;
31734: pixelout<=1'b1;
31735: pixelout<=1'b1;
31736: pixelout<=1'b1;
31737: pixelout<=1'b1;
31738: pixelout<=1'b1;
31739: pixelout<=1'b1;
31740: pixelout<=1'b1;
31741: pixelout<=1'b1;
31742: pixelout<=1'b1;
31743: pixelout<=1'b1;
31744: pixelout<=1'b1;
31745: pixelout<=1'b1;
31746: pixelout<=1'b1;
31747: pixelout<=1'b1;
31748: pixelout<=1'b1;
31749: pixelout<=1'b1;
31750: pixelout<=1'b1;
31751: pixelout<=1'b1;
31752: pixelout<=1'b1;
31753: pixelout<=1'b1;
31754: pixelout<=1'b1;
31755: pixelout<=1'b0;
31756: pixelout<=1'b1;
31757: pixelout<=1'b1;
31758: pixelout<=1'b1;
31759: pixelout<=1'b1;
31760: pixelout<=1'b1;
31761: pixelout<=1'b1;
31762: pixelout<=1'b1;
31763: pixelout<=1'b1;
31764: pixelout<=1'b1;
31765: pixelout<=1'b1;
31766: pixelout<=1'b1;
31767: pixelout<=1'b1;
31768: pixelout<=1'b1;
31769: pixelout<=1'b1;
31770: pixelout<=1'b1;
31771: pixelout<=1'b1;
31772: pixelout<=1'b1;
31773: pixelout<=1'b1;
31774: pixelout<=1'b1;
31775: pixelout<=1'b1;
31776: pixelout<=1'b1;
31777: pixelout<=1'b1;
31778: pixelout<=1'b1;
31779: pixelout<=1'b1;
31780: pixelout<=1'b1;
31781: pixelout<=1'b1;
31782: pixelout<=1'b1;
31783: pixelout<=1'b1;
31784: pixelout<=1'b1;
31785: pixelout<=1'b1;
31786: pixelout<=1'b1;
31787: pixelout<=1'b1;
31788: pixelout<=1'b1;
31789: pixelout<=1'b1;
31790: pixelout<=1'b1;
31791: pixelout<=1'b1;
31792: pixelout<=1'b1;
31793: pixelout<=1'b1;
31794: pixelout<=1'b1;
31795: pixelout<=1'b1;
31796: pixelout<=1'b1;
31797: pixelout<=1'b1;
31798: pixelout<=1'b1;
31799: pixelout<=1'b1;
31800: pixelout<=1'b1;
31801: pixelout<=1'b1;
31802: pixelout<=1'b1;
31803: pixelout<=1'b1;
31804: pixelout<=1'b1;
31805: pixelout<=1'b1;
31806: pixelout<=1'b1;
31807: pixelout<=1'b1;
31808: pixelout<=1'b1;
31809: pixelout<=1'b0;
31810: pixelout<=1'b1;
31811: pixelout<=1'b1;
31812: pixelout<=1'b1;
31813: pixelout<=1'b0;
31814: pixelout<=1'b1;
31815: pixelout<=1'b1;
31816: pixelout<=1'b1;
31817: pixelout<=1'b1;
31818: pixelout<=1'b1;
31819: pixelout<=1'b1;
31820: pixelout<=1'b1;
31821: pixelout<=1'b1;
31822: pixelout<=1'b1;
31823: pixelout<=1'b1;
31824: pixelout<=1'b1;
31825: pixelout<=1'b1;
31826: pixelout<=1'b1;
31827: pixelout<=1'b1;
31828: pixelout<=1'b1;
31829: pixelout<=1'b1;
31830: pixelout<=1'b1;
31831: pixelout<=1'b1;
31832: pixelout<=1'b1;
31833: pixelout<=1'b1;
31834: pixelout<=1'b1;
31835: pixelout<=1'b1;
31836: pixelout<=1'b1;
31837: pixelout<=1'b1;
31838: pixelout<=1'b1;
31839: pixelout<=1'b1;
31840: pixelout<=1'b1;
31841: pixelout<=1'b1;
31842: pixelout<=1'b1;
31843: pixelout<=1'b1;
31844: pixelout<=1'b1;
31845: pixelout<=1'b1;
31846: pixelout<=1'b1;
31847: pixelout<=1'b1;
31848: pixelout<=1'b1;
31849: pixelout<=1'b1;
31850: pixelout<=1'b1;
31851: pixelout<=1'b0;
31852: pixelout<=1'b1;
31853: pixelout<=1'b1;
31854: pixelout<=1'b1;
31855: pixelout<=1'b0;
31856: pixelout<=1'b1;
31857: pixelout<=1'b1;
31858: pixelout<=1'b1;
31859: pixelout<=1'b1;
31860: pixelout<=1'b1;
31861: pixelout<=1'b1;
31862: pixelout<=1'b1;
31863: pixelout<=1'b1;
31864: pixelout<=1'b1;
31865: pixelout<=1'b1;
31866: pixelout<=1'b1;
31867: pixelout<=1'b1;
31868: pixelout<=1'b1;
31869: pixelout<=1'b1;
31870: pixelout<=1'b0;
31871: pixelout<=1'b1;
31872: pixelout<=1'b1;
31873: pixelout<=1'b1;
31874: pixelout<=1'b1;
31875: pixelout<=1'b1;
31876: pixelout<=1'b1;
31877: pixelout<=1'b1;
31878: pixelout<=1'b1;
31879: pixelout<=1'b1;
31880: pixelout<=1'b1;
31881: pixelout<=1'b1;
31882: pixelout<=1'b1;
31883: pixelout<=1'b1;
31884: pixelout<=1'b1;
31885: pixelout<=1'b1;
31886: pixelout<=1'b1;
31887: pixelout<=1'b1;
31888: pixelout<=1'b1;
31889: pixelout<=1'b1;
31890: pixelout<=1'b1;
31891: pixelout<=1'b1;
31892: pixelout<=1'b1;
31893: pixelout<=1'b1;
31894: pixelout<=1'b1;
31895: pixelout<=1'b1;
31896: pixelout<=1'b1;
31897: pixelout<=1'b1;
31898: pixelout<=1'b1;
31899: pixelout<=1'b1;
31900: pixelout<=1'b1;
31901: pixelout<=1'b1;
31902: pixelout<=1'b1;
31903: pixelout<=1'b1;
31904: pixelout<=1'b1;
31905: pixelout<=1'b1;
31906: pixelout<=1'b1;
31907: pixelout<=1'b1;
31908: pixelout<=1'b1;
31909: pixelout<=1'b1;
31910: pixelout<=1'b1;
31911: pixelout<=1'b1;
31912: pixelout<=1'b1;
31913: pixelout<=1'b1;
31914: pixelout<=1'b1;
31915: pixelout<=1'b1;
31916: pixelout<=1'b1;
31917: pixelout<=1'b1;
31918: pixelout<=1'b1;
31919: pixelout<=1'b1;
31920: pixelout<=1'b1;
31921: pixelout<=1'b1;
31922: pixelout<=1'b1;
31923: pixelout<=1'b1;
31924: pixelout<=1'b1;
31925: pixelout<=1'b1;
31926: pixelout<=1'b1;
31927: pixelout<=1'b1;
31928: pixelout<=1'b1;
31929: pixelout<=1'b1;
31930: pixelout<=1'b1;
31931: pixelout<=1'b1;
31932: pixelout<=1'b1;
31933: pixelout<=1'b1;
31934: pixelout<=1'b1;
31935: pixelout<=1'b1;
31936: pixelout<=1'b1;
31937: pixelout<=1'b1;
31938: pixelout<=1'b1;
31939: pixelout<=1'b1;
31940: pixelout<=1'b1;
31941: pixelout<=1'b1;
31942: pixelout<=1'b1;
31943: pixelout<=1'b1;
31944: pixelout<=1'b1;
31945: pixelout<=1'b1;
31946: pixelout<=1'b1;
31947: pixelout<=1'b1;
31948: pixelout<=1'b1;
31949: pixelout<=1'b1;
31950: pixelout<=1'b1;
31951: pixelout<=1'b1;
31952: pixelout<=1'b1;
31953: pixelout<=1'b1;
31954: pixelout<=1'b1;
31955: pixelout<=1'b1;
31956: pixelout<=1'b1;
31957: pixelout<=1'b1;
31958: pixelout<=1'b1;
31959: pixelout<=1'b1;
31960: pixelout<=1'b1;
31961: pixelout<=1'b1;
31962: pixelout<=1'b1;
31963: pixelout<=1'b0;
31964: pixelout<=1'b0;
31965: pixelout<=1'b0;
31966: pixelout<=1'b0;
31967: pixelout<=1'b1;
31968: pixelout<=1'b1;
31969: pixelout<=1'b1;
31970: pixelout<=1'b1;
31971: pixelout<=1'b0;
31972: pixelout<=1'b0;
31973: pixelout<=1'b0;
31974: pixelout<=1'b1;
31975: pixelout<=1'b1;
31976: pixelout<=1'b0;
31977: pixelout<=1'b1;
31978: pixelout<=1'b0;
31979: pixelout<=1'b0;
31980: pixelout<=1'b1;
31981: pixelout<=1'b1;
31982: pixelout<=1'b1;
31983: pixelout<=1'b0;
31984: pixelout<=1'b0;
31985: pixelout<=1'b1;
31986: pixelout<=1'b1;
31987: pixelout<=1'b1;
31988: pixelout<=1'b1;
31989: pixelout<=1'b0;
31990: pixelout<=1'b0;
31991: pixelout<=1'b0;
31992: pixelout<=1'b0;
31993: pixelout<=1'b1;
31994: pixelout<=1'b0;
31995: pixelout<=1'b0;
31996: pixelout<=1'b0;
31997: pixelout<=1'b0;
31998: pixelout<=1'b1;
31999: pixelout<=1'b1;
32000: pixelout<=1'b1;
32001: pixelout<=1'b0;
32002: pixelout<=1'b0;
32003: pixelout<=1'b0;
32004: pixelout<=1'b0;
32005: pixelout<=1'b1;
32006: pixelout<=1'b0;
32007: pixelout<=1'b1;
32008: pixelout<=1'b1;
32009: pixelout<=1'b0;
32010: pixelout<=1'b1;
32011: pixelout<=1'b1;
32012: pixelout<=1'b1;
32013: pixelout<=1'b0;
32014: pixelout<=1'b0;
32015: pixelout<=1'b0;
32016: pixelout<=1'b1;
32017: pixelout<=1'b1;
32018: pixelout<=1'b1;
32019: pixelout<=1'b0;
32020: pixelout<=1'b0;
32021: pixelout<=1'b0;
32022: pixelout<=1'b0;
32023: pixelout<=1'b1;
32024: pixelout<=1'b1;
32025: pixelout<=1'b1;
32026: pixelout<=1'b0;
32027: pixelout<=1'b0;
32028: pixelout<=1'b0;
32029: pixelout<=1'b1;
32030: pixelout<=1'b1;
32031: pixelout<=1'b0;
32032: pixelout<=1'b1;
32033: pixelout<=1'b1;
32034: pixelout<=1'b0;
32035: pixelout<=1'b1;
32036: pixelout<=1'b1;
32037: pixelout<=1'b1;
32038: pixelout<=1'b1;
32039: pixelout<=1'b1;
32040: pixelout<=1'b1;
32041: pixelout<=1'b1;
32042: pixelout<=1'b1;
32043: pixelout<=1'b0;
32044: pixelout<=1'b0;
32045: pixelout<=1'b0;
32046: pixelout<=1'b0;
32047: pixelout<=1'b0;
32048: pixelout<=1'b1;
32049: pixelout<=1'b0;
32050: pixelout<=1'b1;
32051: pixelout<=1'b1;
32052: pixelout<=1'b1;
32053: pixelout<=1'b0;
32054: pixelout<=1'b1;
32055: pixelout<=1'b0;
32056: pixelout<=1'b1;
32057: pixelout<=1'b1;
32058: pixelout<=1'b0;
32059: pixelout<=1'b1;
32060: pixelout<=1'b1;
32061: pixelout<=1'b1;
32062: pixelout<=1'b0;
32063: pixelout<=1'b0;
32064: pixelout<=1'b1;
32065: pixelout<=1'b1;
32066: pixelout<=1'b1;
32067: pixelout<=1'b1;
32068: pixelout<=1'b1;
32069: pixelout<=1'b1;
32070: pixelout<=1'b1;
32071: pixelout<=1'b0;
32072: pixelout<=1'b1;
32073: pixelout<=1'b1;
32074: pixelout<=1'b1;
32075: pixelout<=1'b1;
32076: pixelout<=1'b0;
32077: pixelout<=1'b0;
32078: pixelout<=1'b0;
32079: pixelout<=1'b0;
32080: pixelout<=1'b1;
32081: pixelout<=1'b0;
32082: pixelout<=1'b0;
32083: pixelout<=1'b0;
32084: pixelout<=1'b1;
32085: pixelout<=1'b1;
32086: pixelout<=1'b1;
32087: pixelout<=1'b1;
32088: pixelout<=1'b0;
32089: pixelout<=1'b0;
32090: pixelout<=1'b0;
32091: pixelout<=1'b0;
32092: pixelout<=1'b1;
32093: pixelout<=1'b1;
32094: pixelout<=1'b1;
32095: pixelout<=1'b0;
32096: pixelout<=1'b0;
32097: pixelout<=1'b0;
32098: pixelout<=1'b0;
32099: pixelout<=1'b1;
32100: pixelout<=1'b1;
32101: pixelout<=1'b0;
32102: pixelout<=1'b0;
32103: pixelout<=1'b0;
32104: pixelout<=1'b0;
32105: pixelout<=1'b1;
32106: pixelout<=1'b1;
32107: pixelout<=1'b0;
32108: pixelout<=1'b1;
32109: pixelout<=1'b1;
32110: pixelout<=1'b0;
32111: pixelout<=1'b1;
32112: pixelout<=1'b1;
32113: pixelout<=1'b1;
32114: pixelout<=1'b1;
32115: pixelout<=1'b1;
32116: pixelout<=1'b1;
32117: pixelout<=1'b0;
32118: pixelout<=1'b1;
32119: pixelout<=1'b1;
32120: pixelout<=1'b1;
32121: pixelout<=1'b1;
32122: pixelout<=1'b1;
32123: pixelout<=1'b1;
32124: pixelout<=1'b1;
32125: pixelout<=1'b1;
32126: pixelout<=1'b1;
32127: pixelout<=1'b1;
32128: pixelout<=1'b1;
32129: pixelout<=1'b1;
32130: pixelout<=1'b1;
32131: pixelout<=1'b1;
32132: pixelout<=1'b1;
32133: pixelout<=1'b1;
32134: pixelout<=1'b1;
32135: pixelout<=1'b1;
32136: pixelout<=1'b1;
32137: pixelout<=1'b1;
32138: pixelout<=1'b1;
32139: pixelout<=1'b1;
32140: pixelout<=1'b1;
32141: pixelout<=1'b1;
32142: pixelout<=1'b1;
32143: pixelout<=1'b1;
32144: pixelout<=1'b1;
32145: pixelout<=1'b1;
32146: pixelout<=1'b1;
32147: pixelout<=1'b1;
32148: pixelout<=1'b1;
32149: pixelout<=1'b1;
32150: pixelout<=1'b1;
32151: pixelout<=1'b1;
32152: pixelout<=1'b1;
32153: pixelout<=1'b1;
32154: pixelout<=1'b1;
32155: pixelout<=1'b1;
32156: pixelout<=1'b1;
32157: pixelout<=1'b1;
32158: pixelout<=1'b1;
32159: pixelout<=1'b1;
32160: pixelout<=1'b1;
32161: pixelout<=1'b1;
32162: pixelout<=1'b1;
32163: pixelout<=1'b1;
32164: pixelout<=1'b1;
32165: pixelout<=1'b1;
32166: pixelout<=1'b1;
32167: pixelout<=1'b1;
32168: pixelout<=1'b1;
32169: pixelout<=1'b1;
32170: pixelout<=1'b1;
32171: pixelout<=1'b1;
32172: pixelout<=1'b1;
32173: pixelout<=1'b1;
32174: pixelout<=1'b1;
32175: pixelout<=1'b1;
32176: pixelout<=1'b1;
32177: pixelout<=1'b1;
32178: pixelout<=1'b1;
32179: pixelout<=1'b1;
32180: pixelout<=1'b1;
32181: pixelout<=1'b1;
32182: pixelout<=1'b1;
32183: pixelout<=1'b1;
32184: pixelout<=1'b1;
32185: pixelout<=1'b1;
32186: pixelout<=1'b1;
32187: pixelout<=1'b1;
32188: pixelout<=1'b1;
32189: pixelout<=1'b1;
32190: pixelout<=1'b1;
32191: pixelout<=1'b1;
32192: pixelout<=1'b1;
32193: pixelout<=1'b1;
32194: pixelout<=1'b1;
32195: pixelout<=1'b1;
32196: pixelout<=1'b1;
32197: pixelout<=1'b1;
32198: pixelout<=1'b1;
32199: pixelout<=1'b1;
32200: pixelout<=1'b1;
32201: pixelout<=1'b1;
32202: pixelout<=1'b1;
32203: pixelout<=1'b1;
32204: pixelout<=1'b1;
32205: pixelout<=1'b1;
32206: pixelout<=1'b0;
32207: pixelout<=1'b1;
32208: pixelout<=1'b1;
32209: pixelout<=1'b1;
32210: pixelout<=1'b0;
32211: pixelout<=1'b1;
32212: pixelout<=1'b1;
32213: pixelout<=1'b1;
32214: pixelout<=1'b0;
32215: pixelout<=1'b1;
32216: pixelout<=1'b0;
32217: pixelout<=1'b0;
32218: pixelout<=1'b1;
32219: pixelout<=1'b1;
32220: pixelout<=1'b1;
32221: pixelout<=1'b0;
32222: pixelout<=1'b1;
32223: pixelout<=1'b1;
32224: pixelout<=1'b1;
32225: pixelout<=1'b1;
32226: pixelout<=1'b1;
32227: pixelout<=1'b1;
32228: pixelout<=1'b1;
32229: pixelout<=1'b1;
32230: pixelout<=1'b1;
32231: pixelout<=1'b1;
32232: pixelout<=1'b0;
32233: pixelout<=1'b1;
32234: pixelout<=1'b1;
32235: pixelout<=1'b0;
32236: pixelout<=1'b1;
32237: pixelout<=1'b1;
32238: pixelout<=1'b1;
32239: pixelout<=1'b1;
32240: pixelout<=1'b1;
32241: pixelout<=1'b0;
32242: pixelout<=1'b1;
32243: pixelout<=1'b1;
32244: pixelout<=1'b1;
32245: pixelout<=1'b1;
32246: pixelout<=1'b0;
32247: pixelout<=1'b1;
32248: pixelout<=1'b1;
32249: pixelout<=1'b0;
32250: pixelout<=1'b1;
32251: pixelout<=1'b1;
32252: pixelout<=1'b1;
32253: pixelout<=1'b1;
32254: pixelout<=1'b1;
32255: pixelout<=1'b0;
32256: pixelout<=1'b1;
32257: pixelout<=1'b0;
32258: pixelout<=1'b1;
32259: pixelout<=1'b0;
32260: pixelout<=1'b1;
32261: pixelout<=1'b0;
32262: pixelout<=1'b1;
32263: pixelout<=1'b0;
32264: pixelout<=1'b1;
32265: pixelout<=1'b0;
32266: pixelout<=1'b1;
32267: pixelout<=1'b1;
32268: pixelout<=1'b1;
32269: pixelout<=1'b0;
32270: pixelout<=1'b1;
32271: pixelout<=1'b0;
32272: pixelout<=1'b0;
32273: pixelout<=1'b1;
32274: pixelout<=1'b1;
32275: pixelout<=1'b1;
32276: pixelout<=1'b1;
32277: pixelout<=1'b1;
32278: pixelout<=1'b1;
32279: pixelout<=1'b1;
32280: pixelout<=1'b1;
32281: pixelout<=1'b1;
32282: pixelout<=1'b1;
32283: pixelout<=1'b1;
32284: pixelout<=1'b1;
32285: pixelout<=1'b1;
32286: pixelout<=1'b1;
32287: pixelout<=1'b1;
32288: pixelout<=1'b1;
32289: pixelout<=1'b0;
32290: pixelout<=1'b0;
32291: pixelout<=1'b0;
32292: pixelout<=1'b0;
32293: pixelout<=1'b0;
32294: pixelout<=1'b1;
32295: pixelout<=1'b0;
32296: pixelout<=1'b0;
32297: pixelout<=1'b1;
32298: pixelout<=1'b1;
32299: pixelout<=1'b1;
32300: pixelout<=1'b0;
32301: pixelout<=1'b1;
32302: pixelout<=1'b1;
32303: pixelout<=1'b1;
32304: pixelout<=1'b1;
32305: pixelout<=1'b1;
32306: pixelout<=1'b1;
32307: pixelout<=1'b1;
32308: pixelout<=1'b1;
32309: pixelout<=1'b1;
32310: pixelout<=1'b1;
32311: pixelout<=1'b0;
32312: pixelout<=1'b1;
32313: pixelout<=1'b1;
32314: pixelout<=1'b1;
32315: pixelout<=1'b0;
32316: pixelout<=1'b1;
32317: pixelout<=1'b1;
32318: pixelout<=1'b1;
32319: pixelout<=1'b0;
32320: pixelout<=1'b1;
32321: pixelout<=1'b0;
32322: pixelout<=1'b1;
32323: pixelout<=1'b1;
32324: pixelout<=1'b0;
32325: pixelout<=1'b1;
32326: pixelout<=1'b1;
32327: pixelout<=1'b1;
32328: pixelout<=1'b1;
32329: pixelout<=1'b1;
32330: pixelout<=1'b1;
32331: pixelout<=1'b0;
32332: pixelout<=1'b1;
32333: pixelout<=1'b1;
32334: pixelout<=1'b1;
32335: pixelout<=1'b0;
32336: pixelout<=1'b1;
32337: pixelout<=1'b1;
32338: pixelout<=1'b1;
32339: pixelout<=1'b1;
32340: pixelout<=1'b1;
32341: pixelout<=1'b0;
32342: pixelout<=1'b1;
32343: pixelout<=1'b0;
32344: pixelout<=1'b1;
32345: pixelout<=1'b0;
32346: pixelout<=1'b1;
32347: pixelout<=1'b0;
32348: pixelout<=1'b1;
32349: pixelout<=1'b1;
32350: pixelout<=1'b0;
32351: pixelout<=1'b1;
32352: pixelout<=1'b1;
32353: pixelout<=1'b1;
32354: pixelout<=1'b1;
32355: pixelout<=1'b1;
32356: pixelout<=1'b1;
32357: pixelout<=1'b0;
32358: pixelout<=1'b1;
32359: pixelout<=1'b1;
32360: pixelout<=1'b1;
32361: pixelout<=1'b1;
32362: pixelout<=1'b1;
32363: pixelout<=1'b1;
32364: pixelout<=1'b1;
32365: pixelout<=1'b1;
32366: pixelout<=1'b1;
32367: pixelout<=1'b1;
32368: pixelout<=1'b1;
32369: pixelout<=1'b1;
32370: pixelout<=1'b1;
32371: pixelout<=1'b1;
32372: pixelout<=1'b1;
32373: pixelout<=1'b1;
32374: pixelout<=1'b1;
32375: pixelout<=1'b1;
32376: pixelout<=1'b1;
32377: pixelout<=1'b1;
32378: pixelout<=1'b1;
32379: pixelout<=1'b1;
32380: pixelout<=1'b1;
32381: pixelout<=1'b1;
32382: pixelout<=1'b1;
32383: pixelout<=1'b1;
32384: pixelout<=1'b1;
32385: pixelout<=1'b1;
32386: pixelout<=1'b1;
32387: pixelout<=1'b1;
32388: pixelout<=1'b1;
32389: pixelout<=1'b1;
32390: pixelout<=1'b1;
32391: pixelout<=1'b1;
32392: pixelout<=1'b1;
32393: pixelout<=1'b1;
32394: pixelout<=1'b1;
32395: pixelout<=1'b1;
32396: pixelout<=1'b1;
32397: pixelout<=1'b1;
32398: pixelout<=1'b1;
32399: pixelout<=1'b1;
32400: pixelout<=1'b1;
32401: pixelout<=1'b1;
32402: pixelout<=1'b1;
32403: pixelout<=1'b1;
32404: pixelout<=1'b1;
32405: pixelout<=1'b1;
32406: pixelout<=1'b1;
32407: pixelout<=1'b1;
32408: pixelout<=1'b1;
32409: pixelout<=1'b1;
32410: pixelout<=1'b1;
32411: pixelout<=1'b1;
32412: pixelout<=1'b1;
32413: pixelout<=1'b1;
32414: pixelout<=1'b1;
32415: pixelout<=1'b1;
32416: pixelout<=1'b1;
32417: pixelout<=1'b1;
32418: pixelout<=1'b1;
32419: pixelout<=1'b1;
32420: pixelout<=1'b1;
32421: pixelout<=1'b1;
32422: pixelout<=1'b1;
32423: pixelout<=1'b1;
32424: pixelout<=1'b1;
32425: pixelout<=1'b1;
32426: pixelout<=1'b1;
32427: pixelout<=1'b1;
32428: pixelout<=1'b1;
32429: pixelout<=1'b1;
32430: pixelout<=1'b1;
32431: pixelout<=1'b1;
32432: pixelout<=1'b1;
32433: pixelout<=1'b1;
32434: pixelout<=1'b1;
32435: pixelout<=1'b1;
32436: pixelout<=1'b1;
32437: pixelout<=1'b1;
32438: pixelout<=1'b1;
32439: pixelout<=1'b1;
32440: pixelout<=1'b1;
32441: pixelout<=1'b1;
32442: pixelout<=1'b1;
32443: pixelout<=1'b1;
32444: pixelout<=1'b1;
32445: pixelout<=1'b1;
32446: pixelout<=1'b0;
32447: pixelout<=1'b1;
32448: pixelout<=1'b1;
32449: pixelout<=1'b1;
32450: pixelout<=1'b0;
32451: pixelout<=1'b1;
32452: pixelout<=1'b1;
32453: pixelout<=1'b1;
32454: pixelout<=1'b0;
32455: pixelout<=1'b1;
32456: pixelout<=1'b0;
32457: pixelout<=1'b1;
32458: pixelout<=1'b1;
32459: pixelout<=1'b1;
32460: pixelout<=1'b1;
32461: pixelout<=1'b0;
32462: pixelout<=1'b0;
32463: pixelout<=1'b0;
32464: pixelout<=1'b0;
32465: pixelout<=1'b0;
32466: pixelout<=1'b1;
32467: pixelout<=1'b1;
32468: pixelout<=1'b1;
32469: pixelout<=1'b1;
32470: pixelout<=1'b1;
32471: pixelout<=1'b1;
32472: pixelout<=1'b0;
32473: pixelout<=1'b1;
32474: pixelout<=1'b1;
32475: pixelout<=1'b0;
32476: pixelout<=1'b1;
32477: pixelout<=1'b1;
32478: pixelout<=1'b1;
32479: pixelout<=1'b1;
32480: pixelout<=1'b1;
32481: pixelout<=1'b1;
32482: pixelout<=1'b0;
32483: pixelout<=1'b0;
32484: pixelout<=1'b1;
32485: pixelout<=1'b1;
32486: pixelout<=1'b0;
32487: pixelout<=1'b1;
32488: pixelout<=1'b1;
32489: pixelout<=1'b0;
32490: pixelout<=1'b1;
32491: pixelout<=1'b1;
32492: pixelout<=1'b1;
32493: pixelout<=1'b1;
32494: pixelout<=1'b1;
32495: pixelout<=1'b0;
32496: pixelout<=1'b1;
32497: pixelout<=1'b0;
32498: pixelout<=1'b1;
32499: pixelout<=1'b0;
32500: pixelout<=1'b1;
32501: pixelout<=1'b0;
32502: pixelout<=1'b1;
32503: pixelout<=1'b0;
32504: pixelout<=1'b1;
32505: pixelout<=1'b0;
32506: pixelout<=1'b0;
32507: pixelout<=1'b0;
32508: pixelout<=1'b0;
32509: pixelout<=1'b0;
32510: pixelout<=1'b1;
32511: pixelout<=1'b0;
32512: pixelout<=1'b1;
32513: pixelout<=1'b1;
32514: pixelout<=1'b1;
32515: pixelout<=1'b1;
32516: pixelout<=1'b1;
32517: pixelout<=1'b1;
32518: pixelout<=1'b1;
32519: pixelout<=1'b1;
32520: pixelout<=1'b1;
32521: pixelout<=1'b1;
32522: pixelout<=1'b1;
32523: pixelout<=1'b1;
32524: pixelout<=1'b1;
32525: pixelout<=1'b1;
32526: pixelout<=1'b1;
32527: pixelout<=1'b1;
32528: pixelout<=1'b1;
32529: pixelout<=1'b0;
32530: pixelout<=1'b1;
32531: pixelout<=1'b1;
32532: pixelout<=1'b1;
32533: pixelout<=1'b0;
32534: pixelout<=1'b1;
32535: pixelout<=1'b0;
32536: pixelout<=1'b1;
32537: pixelout<=1'b1;
32538: pixelout<=1'b1;
32539: pixelout<=1'b1;
32540: pixelout<=1'b0;
32541: pixelout<=1'b1;
32542: pixelout<=1'b1;
32543: pixelout<=1'b1;
32544: pixelout<=1'b1;
32545: pixelout<=1'b1;
32546: pixelout<=1'b1;
32547: pixelout<=1'b1;
32548: pixelout<=1'b1;
32549: pixelout<=1'b1;
32550: pixelout<=1'b1;
32551: pixelout<=1'b0;
32552: pixelout<=1'b1;
32553: pixelout<=1'b1;
32554: pixelout<=1'b1;
32555: pixelout<=1'b0;
32556: pixelout<=1'b1;
32557: pixelout<=1'b1;
32558: pixelout<=1'b1;
32559: pixelout<=1'b0;
32560: pixelout<=1'b1;
32561: pixelout<=1'b0;
32562: pixelout<=1'b1;
32563: pixelout<=1'b1;
32564: pixelout<=1'b0;
32565: pixelout<=1'b1;
32566: pixelout<=1'b1;
32567: pixelout<=1'b1;
32568: pixelout<=1'b1;
32569: pixelout<=1'b1;
32570: pixelout<=1'b1;
32571: pixelout<=1'b0;
32572: pixelout<=1'b1;
32573: pixelout<=1'b1;
32574: pixelout<=1'b1;
32575: pixelout<=1'b0;
32576: pixelout<=1'b1;
32577: pixelout<=1'b1;
32578: pixelout<=1'b1;
32579: pixelout<=1'b1;
32580: pixelout<=1'b1;
32581: pixelout<=1'b0;
32582: pixelout<=1'b1;
32583: pixelout<=1'b0;
32584: pixelout<=1'b1;
32585: pixelout<=1'b0;
32586: pixelout<=1'b1;
32587: pixelout<=1'b0;
32588: pixelout<=1'b1;
32589: pixelout<=1'b1;
32590: pixelout<=1'b0;
32591: pixelout<=1'b1;
32592: pixelout<=1'b1;
32593: pixelout<=1'b1;
32594: pixelout<=1'b1;
32595: pixelout<=1'b1;
32596: pixelout<=1'b1;
32597: pixelout<=1'b0;
32598: pixelout<=1'b1;
32599: pixelout<=1'b1;
32600: pixelout<=1'b1;
32601: pixelout<=1'b1;
32602: pixelout<=1'b1;
32603: pixelout<=1'b1;
32604: pixelout<=1'b1;
32605: pixelout<=1'b1;
32606: pixelout<=1'b1;
32607: pixelout<=1'b1;
32608: pixelout<=1'b1;
32609: pixelout<=1'b1;
32610: pixelout<=1'b1;
32611: pixelout<=1'b1;
32612: pixelout<=1'b1;
32613: pixelout<=1'b1;
32614: pixelout<=1'b1;
32615: pixelout<=1'b1;
32616: pixelout<=1'b1;
32617: pixelout<=1'b1;
32618: pixelout<=1'b1;
32619: pixelout<=1'b1;
32620: pixelout<=1'b1;
32621: pixelout<=1'b1;
32622: pixelout<=1'b1;
32623: pixelout<=1'b1;
32624: pixelout<=1'b1;
32625: pixelout<=1'b1;
32626: pixelout<=1'b1;
32627: pixelout<=1'b1;
32628: pixelout<=1'b1;
32629: pixelout<=1'b1;
32630: pixelout<=1'b1;
32631: pixelout<=1'b1;
32632: pixelout<=1'b1;
32633: pixelout<=1'b1;
32634: pixelout<=1'b1;
32635: pixelout<=1'b1;
32636: pixelout<=1'b1;
32637: pixelout<=1'b1;
32638: pixelout<=1'b1;
32639: pixelout<=1'b1;
32640: pixelout<=1'b1;
32641: pixelout<=1'b1;
32642: pixelout<=1'b1;
32643: pixelout<=1'b1;
32644: pixelout<=1'b1;
32645: pixelout<=1'b1;
32646: pixelout<=1'b1;
32647: pixelout<=1'b1;
32648: pixelout<=1'b1;
32649: pixelout<=1'b1;
32650: pixelout<=1'b1;
32651: pixelout<=1'b1;
32652: pixelout<=1'b1;
32653: pixelout<=1'b1;
32654: pixelout<=1'b1;
32655: pixelout<=1'b1;
32656: pixelout<=1'b1;
32657: pixelout<=1'b1;
32658: pixelout<=1'b1;
32659: pixelout<=1'b1;
32660: pixelout<=1'b1;
32661: pixelout<=1'b1;
32662: pixelout<=1'b1;
32663: pixelout<=1'b1;
32664: pixelout<=1'b1;
32665: pixelout<=1'b1;
32666: pixelout<=1'b1;
32667: pixelout<=1'b1;
32668: pixelout<=1'b1;
32669: pixelout<=1'b1;
32670: pixelout<=1'b1;
32671: pixelout<=1'b1;
32672: pixelout<=1'b1;
32673: pixelout<=1'b1;
32674: pixelout<=1'b1;
32675: pixelout<=1'b1;
32676: pixelout<=1'b1;
32677: pixelout<=1'b1;
32678: pixelout<=1'b1;
32679: pixelout<=1'b1;
32680: pixelout<=1'b1;
32681: pixelout<=1'b1;
32682: pixelout<=1'b1;
32683: pixelout<=1'b1;
32684: pixelout<=1'b1;
32685: pixelout<=1'b0;
32686: pixelout<=1'b0;
32687: pixelout<=1'b1;
32688: pixelout<=1'b1;
32689: pixelout<=1'b1;
32690: pixelout<=1'b0;
32691: pixelout<=1'b1;
32692: pixelout<=1'b1;
32693: pixelout<=1'b1;
32694: pixelout<=1'b0;
32695: pixelout<=1'b1;
32696: pixelout<=1'b0;
32697: pixelout<=1'b1;
32698: pixelout<=1'b1;
32699: pixelout<=1'b1;
32700: pixelout<=1'b1;
32701: pixelout<=1'b0;
32702: pixelout<=1'b1;
32703: pixelout<=1'b1;
32704: pixelout<=1'b1;
32705: pixelout<=1'b1;
32706: pixelout<=1'b1;
32707: pixelout<=1'b1;
32708: pixelout<=1'b1;
32709: pixelout<=1'b1;
32710: pixelout<=1'b1;
32711: pixelout<=1'b0;
32712: pixelout<=1'b0;
32713: pixelout<=1'b1;
32714: pixelout<=1'b1;
32715: pixelout<=1'b0;
32716: pixelout<=1'b1;
32717: pixelout<=1'b1;
32718: pixelout<=1'b1;
32719: pixelout<=1'b1;
32720: pixelout<=1'b1;
32721: pixelout<=1'b1;
32722: pixelout<=1'b1;
32723: pixelout<=1'b1;
32724: pixelout<=1'b0;
32725: pixelout<=1'b1;
32726: pixelout<=1'b0;
32727: pixelout<=1'b1;
32728: pixelout<=1'b1;
32729: pixelout<=1'b0;
32730: pixelout<=1'b1;
32731: pixelout<=1'b1;
32732: pixelout<=1'b1;
32733: pixelout<=1'b1;
32734: pixelout<=1'b1;
32735: pixelout<=1'b0;
32736: pixelout<=1'b1;
32737: pixelout<=1'b0;
32738: pixelout<=1'b1;
32739: pixelout<=1'b0;
32740: pixelout<=1'b1;
32741: pixelout<=1'b0;
32742: pixelout<=1'b1;
32743: pixelout<=1'b0;
32744: pixelout<=1'b1;
32745: pixelout<=1'b0;
32746: pixelout<=1'b1;
32747: pixelout<=1'b1;
32748: pixelout<=1'b1;
32749: pixelout<=1'b1;
32750: pixelout<=1'b1;
32751: pixelout<=1'b0;
32752: pixelout<=1'b1;
32753: pixelout<=1'b1;
32754: pixelout<=1'b1;
32755: pixelout<=1'b1;
32756: pixelout<=1'b1;
32757: pixelout<=1'b1;
32758: pixelout<=1'b1;
32759: pixelout<=1'b1;
32760: pixelout<=1'b1;
32761: pixelout<=1'b1;
32762: pixelout<=1'b1;
32763: pixelout<=1'b1;
32764: pixelout<=1'b1;
32765: pixelout<=1'b1;
32766: pixelout<=1'b1;
32767: pixelout<=1'b1;
32768: pixelout<=1'b1;
32769: pixelout<=1'b0;
32770: pixelout<=1'b1;
32771: pixelout<=1'b1;
32772: pixelout<=1'b1;
32773: pixelout<=1'b0;
32774: pixelout<=1'b1;
32775: pixelout<=1'b0;
32776: pixelout<=1'b1;
32777: pixelout<=1'b1;
32778: pixelout<=1'b1;
32779: pixelout<=1'b1;
32780: pixelout<=1'b0;
32781: pixelout<=1'b1;
32782: pixelout<=1'b1;
32783: pixelout<=1'b1;
32784: pixelout<=1'b1;
32785: pixelout<=1'b1;
32786: pixelout<=1'b1;
32787: pixelout<=1'b1;
32788: pixelout<=1'b1;
32789: pixelout<=1'b1;
32790: pixelout<=1'b1;
32791: pixelout<=1'b0;
32792: pixelout<=1'b1;
32793: pixelout<=1'b1;
32794: pixelout<=1'b1;
32795: pixelout<=1'b0;
32796: pixelout<=1'b1;
32797: pixelout<=1'b1;
32798: pixelout<=1'b0;
32799: pixelout<=1'b0;
32800: pixelout<=1'b1;
32801: pixelout<=1'b0;
32802: pixelout<=1'b1;
32803: pixelout<=1'b1;
32804: pixelout<=1'b0;
32805: pixelout<=1'b1;
32806: pixelout<=1'b1;
32807: pixelout<=1'b1;
32808: pixelout<=1'b1;
32809: pixelout<=1'b1;
32810: pixelout<=1'b1;
32811: pixelout<=1'b0;
32812: pixelout<=1'b1;
32813: pixelout<=1'b1;
32814: pixelout<=1'b1;
32815: pixelout<=1'b0;
32816: pixelout<=1'b1;
32817: pixelout<=1'b1;
32818: pixelout<=1'b1;
32819: pixelout<=1'b1;
32820: pixelout<=1'b1;
32821: pixelout<=1'b0;
32822: pixelout<=1'b1;
32823: pixelout<=1'b0;
32824: pixelout<=1'b1;
32825: pixelout<=1'b0;
32826: pixelout<=1'b1;
32827: pixelout<=1'b0;
32828: pixelout<=1'b1;
32829: pixelout<=1'b1;
32830: pixelout<=1'b0;
32831: pixelout<=1'b1;
32832: pixelout<=1'b1;
32833: pixelout<=1'b1;
32834: pixelout<=1'b1;
32835: pixelout<=1'b1;
32836: pixelout<=1'b1;
32837: pixelout<=1'b0;
32838: pixelout<=1'b1;
32839: pixelout<=1'b1;
32840: pixelout<=1'b1;
32841: pixelout<=1'b1;
32842: pixelout<=1'b1;
32843: pixelout<=1'b1;
32844: pixelout<=1'b1;
32845: pixelout<=1'b1;
32846: pixelout<=1'b1;
32847: pixelout<=1'b1;
32848: pixelout<=1'b1;
32849: pixelout<=1'b1;
32850: pixelout<=1'b1;
32851: pixelout<=1'b1;
32852: pixelout<=1'b1;
32853: pixelout<=1'b1;
32854: pixelout<=1'b1;
32855: pixelout<=1'b1;
32856: pixelout<=1'b1;
32857: pixelout<=1'b1;
32858: pixelout<=1'b1;
32859: pixelout<=1'b1;
32860: pixelout<=1'b1;
32861: pixelout<=1'b1;
32862: pixelout<=1'b1;
32863: pixelout<=1'b1;
32864: pixelout<=1'b1;
32865: pixelout<=1'b1;
32866: pixelout<=1'b1;
32867: pixelout<=1'b1;
32868: pixelout<=1'b1;
32869: pixelout<=1'b1;
32870: pixelout<=1'b1;
32871: pixelout<=1'b1;
32872: pixelout<=1'b1;
32873: pixelout<=1'b1;
32874: pixelout<=1'b1;
32875: pixelout<=1'b1;
32876: pixelout<=1'b1;
32877: pixelout<=1'b1;
32878: pixelout<=1'b1;
32879: pixelout<=1'b1;
32880: pixelout<=1'b1;
32881: pixelout<=1'b1;
32882: pixelout<=1'b1;
32883: pixelout<=1'b1;
32884: pixelout<=1'b1;
32885: pixelout<=1'b1;
32886: pixelout<=1'b1;
32887: pixelout<=1'b1;
32888: pixelout<=1'b1;
32889: pixelout<=1'b1;
32890: pixelout<=1'b1;
32891: pixelout<=1'b1;
32892: pixelout<=1'b1;
32893: pixelout<=1'b1;
32894: pixelout<=1'b1;
32895: pixelout<=1'b1;
32896: pixelout<=1'b1;
32897: pixelout<=1'b1;
32898: pixelout<=1'b1;
32899: pixelout<=1'b1;
32900: pixelout<=1'b1;
32901: pixelout<=1'b1;
32902: pixelout<=1'b1;
32903: pixelout<=1'b1;
32904: pixelout<=1'b1;
32905: pixelout<=1'b1;
32906: pixelout<=1'b1;
32907: pixelout<=1'b1;
32908: pixelout<=1'b1;
32909: pixelout<=1'b1;
32910: pixelout<=1'b1;
32911: pixelout<=1'b1;
32912: pixelout<=1'b1;
32913: pixelout<=1'b1;
32914: pixelout<=1'b1;
32915: pixelout<=1'b1;
32916: pixelout<=1'b1;
32917: pixelout<=1'b1;
32918: pixelout<=1'b1;
32919: pixelout<=1'b1;
32920: pixelout<=1'b1;
32921: pixelout<=1'b1;
32922: pixelout<=1'b1;
32923: pixelout<=1'b0;
32924: pixelout<=1'b0;
32925: pixelout<=1'b1;
32926: pixelout<=1'b0;
32927: pixelout<=1'b1;
32928: pixelout<=1'b1;
32929: pixelout<=1'b1;
32930: pixelout<=1'b1;
32931: pixelout<=1'b0;
32932: pixelout<=1'b0;
32933: pixelout<=1'b0;
32934: pixelout<=1'b0;
32935: pixelout<=1'b1;
32936: pixelout<=1'b0;
32937: pixelout<=1'b1;
32938: pixelout<=1'b1;
32939: pixelout<=1'b1;
32940: pixelout<=1'b1;
32941: pixelout<=1'b1;
32942: pixelout<=1'b0;
32943: pixelout<=1'b0;
32944: pixelout<=1'b0;
32945: pixelout<=1'b0;
32946: pixelout<=1'b1;
32947: pixelout<=1'b1;
32948: pixelout<=1'b1;
32949: pixelout<=1'b0;
32950: pixelout<=1'b0;
32951: pixelout<=1'b1;
32952: pixelout<=1'b0;
32953: pixelout<=1'b1;
32954: pixelout<=1'b1;
32955: pixelout<=1'b0;
32956: pixelout<=1'b0;
32957: pixelout<=1'b0;
32958: pixelout<=1'b1;
32959: pixelout<=1'b1;
32960: pixelout<=1'b1;
32961: pixelout<=1'b0;
32962: pixelout<=1'b0;
32963: pixelout<=1'b0;
32964: pixelout<=1'b0;
32965: pixelout<=1'b1;
32966: pixelout<=1'b1;
32967: pixelout<=1'b0;
32968: pixelout<=1'b0;
32969: pixelout<=1'b1;
32970: pixelout<=1'b1;
32971: pixelout<=1'b1;
32972: pixelout<=1'b1;
32973: pixelout<=1'b1;
32974: pixelout<=1'b1;
32975: pixelout<=1'b0;
32976: pixelout<=1'b1;
32977: pixelout<=1'b0;
32978: pixelout<=1'b1;
32979: pixelout<=1'b0;
32980: pixelout<=1'b1;
32981: pixelout<=1'b0;
32982: pixelout<=1'b1;
32983: pixelout<=1'b0;
32984: pixelout<=1'b1;
32985: pixelout<=1'b1;
32986: pixelout<=1'b0;
32987: pixelout<=1'b0;
32988: pixelout<=1'b0;
32989: pixelout<=1'b0;
32990: pixelout<=1'b1;
32991: pixelout<=1'b0;
32992: pixelout<=1'b1;
32993: pixelout<=1'b1;
32994: pixelout<=1'b1;
32995: pixelout<=1'b1;
32996: pixelout<=1'b1;
32997: pixelout<=1'b1;
32998: pixelout<=1'b1;
32999: pixelout<=1'b1;
33000: pixelout<=1'b1;
33001: pixelout<=1'b1;
33002: pixelout<=1'b1;
33003: pixelout<=1'b1;
33004: pixelout<=1'b1;
33005: pixelout<=1'b1;
33006: pixelout<=1'b1;
33007: pixelout<=1'b1;
33008: pixelout<=1'b1;
33009: pixelout<=1'b0;
33010: pixelout<=1'b1;
33011: pixelout<=1'b1;
33012: pixelout<=1'b1;
33013: pixelout<=1'b0;
33014: pixelout<=1'b1;
33015: pixelout<=1'b0;
33016: pixelout<=1'b1;
33017: pixelout<=1'b1;
33018: pixelout<=1'b1;
33019: pixelout<=1'b1;
33020: pixelout<=1'b1;
33021: pixelout<=1'b0;
33022: pixelout<=1'b0;
33023: pixelout<=1'b0;
33024: pixelout<=1'b1;
33025: pixelout<=1'b1;
33026: pixelout<=1'b1;
33027: pixelout<=1'b1;
33028: pixelout<=1'b0;
33029: pixelout<=1'b0;
33030: pixelout<=1'b0;
33031: pixelout<=1'b0;
33032: pixelout<=1'b1;
33033: pixelout<=1'b1;
33034: pixelout<=1'b1;
33035: pixelout<=1'b1;
33036: pixelout<=1'b0;
33037: pixelout<=1'b0;
33038: pixelout<=1'b1;
33039: pixelout<=1'b0;
33040: pixelout<=1'b1;
33041: pixelout<=1'b0;
33042: pixelout<=1'b1;
33043: pixelout<=1'b1;
33044: pixelout<=1'b0;
33045: pixelout<=1'b1;
33046: pixelout<=1'b1;
33047: pixelout<=1'b1;
33048: pixelout<=1'b0;
33049: pixelout<=1'b0;
33050: pixelout<=1'b0;
33051: pixelout<=1'b0;
33052: pixelout<=1'b1;
33053: pixelout<=1'b1;
33054: pixelout<=1'b1;
33055: pixelout<=1'b0;
33056: pixelout<=1'b0;
33057: pixelout<=1'b0;
33058: pixelout<=1'b0;
33059: pixelout<=1'b0;
33060: pixelout<=1'b1;
33061: pixelout<=1'b0;
33062: pixelout<=1'b1;
33063: pixelout<=1'b0;
33064: pixelout<=1'b1;
33065: pixelout<=1'b0;
33066: pixelout<=1'b1;
33067: pixelout<=1'b0;
33068: pixelout<=1'b1;
33069: pixelout<=1'b1;
33070: pixelout<=1'b0;
33071: pixelout<=1'b1;
33072: pixelout<=1'b1;
33073: pixelout<=1'b1;
33074: pixelout<=1'b0;
33075: pixelout<=1'b0;
33076: pixelout<=1'b0;
33077: pixelout<=1'b0;
33078: pixelout<=1'b1;
33079: pixelout<=1'b1;
33080: pixelout<=1'b1;
33081: pixelout<=1'b1;
33082: pixelout<=1'b1;
33083: pixelout<=1'b1;
33084: pixelout<=1'b1;
33085: pixelout<=1'b1;
33086: pixelout<=1'b1;
33087: pixelout<=1'b1;
33088: pixelout<=1'b1;
33089: pixelout<=1'b1;
33090: pixelout<=1'b1;
33091: pixelout<=1'b1;
33092: pixelout<=1'b1;
33093: pixelout<=1'b1;
33094: pixelout<=1'b1;
33095: pixelout<=1'b1;
33096: pixelout<=1'b1;
33097: pixelout<=1'b1;
33098: pixelout<=1'b1;
33099: pixelout<=1'b1;
33100: pixelout<=1'b1;
33101: pixelout<=1'b1;
33102: pixelout<=1'b1;
33103: pixelout<=1'b1;
33104: pixelout<=1'b1;
33105: pixelout<=1'b1;
33106: pixelout<=1'b1;
33107: pixelout<=1'b1;
33108: pixelout<=1'b1;
33109: pixelout<=1'b1;
33110: pixelout<=1'b1;
33111: pixelout<=1'b1;
33112: pixelout<=1'b1;
33113: pixelout<=1'b1;
33114: pixelout<=1'b1;
33115: pixelout<=1'b1;
33116: pixelout<=1'b1;
33117: pixelout<=1'b1;
33118: pixelout<=1'b1;
33119: pixelout<=1'b1;
33120: pixelout<=1'b1;
33121: pixelout<=1'b1;
33122: pixelout<=1'b1;
33123: pixelout<=1'b1;
33124: pixelout<=1'b1;
33125: pixelout<=1'b1;
33126: pixelout<=1'b1;
33127: pixelout<=1'b1;
33128: pixelout<=1'b1;
33129: pixelout<=1'b1;
33130: pixelout<=1'b1;
33131: pixelout<=1'b1;
33132: pixelout<=1'b1;
33133: pixelout<=1'b1;
33134: pixelout<=1'b1;
33135: pixelout<=1'b1;
33136: pixelout<=1'b1;
33137: pixelout<=1'b1;
33138: pixelout<=1'b1;
33139: pixelout<=1'b1;
33140: pixelout<=1'b1;
33141: pixelout<=1'b1;
33142: pixelout<=1'b1;
33143: pixelout<=1'b1;
33144: pixelout<=1'b1;
33145: pixelout<=1'b1;
33146: pixelout<=1'b1;
33147: pixelout<=1'b1;
33148: pixelout<=1'b1;
33149: pixelout<=1'b1;
33150: pixelout<=1'b1;
33151: pixelout<=1'b1;
33152: pixelout<=1'b1;
33153: pixelout<=1'b1;
33154: pixelout<=1'b1;
33155: pixelout<=1'b1;
33156: pixelout<=1'b1;
33157: pixelout<=1'b1;
33158: pixelout<=1'b1;
33159: pixelout<=1'b1;
33160: pixelout<=1'b1;
33161: pixelout<=1'b1;
33162: pixelout<=1'b1;
33163: pixelout<=1'b1;
33164: pixelout<=1'b1;
33165: pixelout<=1'b1;
33166: pixelout<=1'b1;
33167: pixelout<=1'b1;
33168: pixelout<=1'b1;
33169: pixelout<=1'b1;
33170: pixelout<=1'b1;
33171: pixelout<=1'b1;
33172: pixelout<=1'b1;
33173: pixelout<=1'b1;
33174: pixelout<=1'b0;
33175: pixelout<=1'b1;
33176: pixelout<=1'b1;
33177: pixelout<=1'b1;
33178: pixelout<=1'b1;
33179: pixelout<=1'b1;
33180: pixelout<=1'b1;
33181: pixelout<=1'b1;
33182: pixelout<=1'b1;
33183: pixelout<=1'b1;
33184: pixelout<=1'b1;
33185: pixelout<=1'b1;
33186: pixelout<=1'b1;
33187: pixelout<=1'b1;
33188: pixelout<=1'b1;
33189: pixelout<=1'b1;
33190: pixelout<=1'b1;
33191: pixelout<=1'b1;
33192: pixelout<=1'b1;
33193: pixelout<=1'b1;
33194: pixelout<=1'b1;
33195: pixelout<=1'b1;
33196: pixelout<=1'b1;
33197: pixelout<=1'b1;
33198: pixelout<=1'b1;
33199: pixelout<=1'b1;
33200: pixelout<=1'b1;
33201: pixelout<=1'b1;
33202: pixelout<=1'b1;
33203: pixelout<=1'b1;
33204: pixelout<=1'b1;
33205: pixelout<=1'b1;
33206: pixelout<=1'b1;
33207: pixelout<=1'b1;
33208: pixelout<=1'b1;
33209: pixelout<=1'b1;
33210: pixelout<=1'b1;
33211: pixelout<=1'b1;
33212: pixelout<=1'b1;
33213: pixelout<=1'b1;
33214: pixelout<=1'b1;
33215: pixelout<=1'b1;
33216: pixelout<=1'b1;
33217: pixelout<=1'b1;
33218: pixelout<=1'b1;
33219: pixelout<=1'b1;
33220: pixelout<=1'b1;
33221: pixelout<=1'b1;
33222: pixelout<=1'b1;
33223: pixelout<=1'b1;
33224: pixelout<=1'b1;
33225: pixelout<=1'b1;
33226: pixelout<=1'b1;
33227: pixelout<=1'b1;
33228: pixelout<=1'b1;
33229: pixelout<=1'b1;
33230: pixelout<=1'b1;
33231: pixelout<=1'b1;
33232: pixelout<=1'b1;
33233: pixelout<=1'b1;
33234: pixelout<=1'b1;
33235: pixelout<=1'b1;
33236: pixelout<=1'b1;
33237: pixelout<=1'b1;
33238: pixelout<=1'b1;
33239: pixelout<=1'b1;
33240: pixelout<=1'b1;
33241: pixelout<=1'b1;
33242: pixelout<=1'b1;
33243: pixelout<=1'b1;
33244: pixelout<=1'b1;
33245: pixelout<=1'b1;
33246: pixelout<=1'b1;
33247: pixelout<=1'b1;
33248: pixelout<=1'b1;
33249: pixelout<=1'b1;
33250: pixelout<=1'b1;
33251: pixelout<=1'b1;
33252: pixelout<=1'b1;
33253: pixelout<=1'b1;
33254: pixelout<=1'b1;
33255: pixelout<=1'b1;
33256: pixelout<=1'b1;
33257: pixelout<=1'b1;
33258: pixelout<=1'b1;
33259: pixelout<=1'b1;
33260: pixelout<=1'b1;
33261: pixelout<=1'b1;
33262: pixelout<=1'b1;
33263: pixelout<=1'b1;
33264: pixelout<=1'b1;
33265: pixelout<=1'b1;
33266: pixelout<=1'b1;
33267: pixelout<=1'b1;
33268: pixelout<=1'b1;
33269: pixelout<=1'b1;
33270: pixelout<=1'b1;
33271: pixelout<=1'b0;
33272: pixelout<=1'b1;
33273: pixelout<=1'b1;
33274: pixelout<=1'b1;
33275: pixelout<=1'b1;
33276: pixelout<=1'b1;
33277: pixelout<=1'b1;
33278: pixelout<=1'b1;
33279: pixelout<=1'b1;
33280: pixelout<=1'b1;
33281: pixelout<=1'b1;
33282: pixelout<=1'b1;
33283: pixelout<=1'b1;
33284: pixelout<=1'b1;
33285: pixelout<=1'b1;
33286: pixelout<=1'b1;
33287: pixelout<=1'b1;
33288: pixelout<=1'b1;
33289: pixelout<=1'b1;
33290: pixelout<=1'b1;
33291: pixelout<=1'b1;
33292: pixelout<=1'b1;
33293: pixelout<=1'b1;
33294: pixelout<=1'b1;
33295: pixelout<=1'b1;
33296: pixelout<=1'b1;
33297: pixelout<=1'b1;
33298: pixelout<=1'b1;
33299: pixelout<=1'b1;
33300: pixelout<=1'b1;
33301: pixelout<=1'b1;
33302: pixelout<=1'b1;
33303: pixelout<=1'b1;
33304: pixelout<=1'b1;
33305: pixelout<=1'b1;
33306: pixelout<=1'b1;
33307: pixelout<=1'b1;
33308: pixelout<=1'b1;
33309: pixelout<=1'b1;
33310: pixelout<=1'b1;
33311: pixelout<=1'b1;
33312: pixelout<=1'b1;
33313: pixelout<=1'b1;
33314: pixelout<=1'b1;
33315: pixelout<=1'b1;
33316: pixelout<=1'b1;
33317: pixelout<=1'b0;
33318: pixelout<=1'b1;
33319: pixelout<=1'b1;
33320: pixelout<=1'b1;
33321: pixelout<=1'b1;
33322: pixelout<=1'b1;
33323: pixelout<=1'b1;
33324: pixelout<=1'b1;
33325: pixelout<=1'b1;
33326: pixelout<=1'b1;
33327: pixelout<=1'b1;
33328: pixelout<=1'b1;
33329: pixelout<=1'b1;
33330: pixelout<=1'b1;
33331: pixelout<=1'b1;
33332: pixelout<=1'b1;
33333: pixelout<=1'b1;
33334: pixelout<=1'b1;
33335: pixelout<=1'b1;
33336: pixelout<=1'b1;
33337: pixelout<=1'b1;
33338: pixelout<=1'b1;
33339: pixelout<=1'b1;
33340: pixelout<=1'b1;
33341: pixelout<=1'b1;
33342: pixelout<=1'b1;
33343: pixelout<=1'b1;
33344: pixelout<=1'b1;
33345: pixelout<=1'b1;
33346: pixelout<=1'b1;
33347: pixelout<=1'b1;
33348: pixelout<=1'b1;
33349: pixelout<=1'b1;
33350: pixelout<=1'b1;
33351: pixelout<=1'b1;
33352: pixelout<=1'b1;
33353: pixelout<=1'b1;
33354: pixelout<=1'b1;
33355: pixelout<=1'b1;
33356: pixelout<=1'b1;
33357: pixelout<=1'b1;
33358: pixelout<=1'b1;
33359: pixelout<=1'b1;
33360: pixelout<=1'b1;
33361: pixelout<=1'b1;
33362: pixelout<=1'b1;
33363: pixelout<=1'b1;
33364: pixelout<=1'b1;
33365: pixelout<=1'b1;
33366: pixelout<=1'b1;
33367: pixelout<=1'b1;
33368: pixelout<=1'b1;
33369: pixelout<=1'b1;
33370: pixelout<=1'b1;
33371: pixelout<=1'b1;
33372: pixelout<=1'b1;
33373: pixelout<=1'b1;
33374: pixelout<=1'b1;
33375: pixelout<=1'b1;
33376: pixelout<=1'b1;
33377: pixelout<=1'b1;
33378: pixelout<=1'b1;
33379: pixelout<=1'b1;
33380: pixelout<=1'b1;
33381: pixelout<=1'b1;
33382: pixelout<=1'b1;
33383: pixelout<=1'b1;
33384: pixelout<=1'b1;
33385: pixelout<=1'b1;
33386: pixelout<=1'b1;
33387: pixelout<=1'b1;
33388: pixelout<=1'b1;
33389: pixelout<=1'b1;
33390: pixelout<=1'b1;
33391: pixelout<=1'b1;
33392: pixelout<=1'b1;
33393: pixelout<=1'b1;
33394: pixelout<=1'b1;
33395: pixelout<=1'b1;
33396: pixelout<=1'b1;
33397: pixelout<=1'b1;
33398: pixelout<=1'b1;
33399: pixelout<=1'b1;
33400: pixelout<=1'b1;
33401: pixelout<=1'b1;
33402: pixelout<=1'b1;
33403: pixelout<=1'b1;
33404: pixelout<=1'b1;
33405: pixelout<=1'b1;
33406: pixelout<=1'b1;
33407: pixelout<=1'b1;
33408: pixelout<=1'b1;
33409: pixelout<=1'b1;
33410: pixelout<=1'b1;
33411: pixelout<=1'b0;
33412: pixelout<=1'b0;
33413: pixelout<=1'b0;
33414: pixelout<=1'b1;
33415: pixelout<=1'b1;
33416: pixelout<=1'b1;
33417: pixelout<=1'b1;
33418: pixelout<=1'b1;
33419: pixelout<=1'b1;
33420: pixelout<=1'b1;
33421: pixelout<=1'b1;
33422: pixelout<=1'b1;
33423: pixelout<=1'b1;
33424: pixelout<=1'b1;
33425: pixelout<=1'b1;
33426: pixelout<=1'b1;
33427: pixelout<=1'b1;
33428: pixelout<=1'b1;
33429: pixelout<=1'b1;
33430: pixelout<=1'b1;
33431: pixelout<=1'b1;
33432: pixelout<=1'b1;
33433: pixelout<=1'b1;
33434: pixelout<=1'b1;
33435: pixelout<=1'b1;
33436: pixelout<=1'b1;
33437: pixelout<=1'b1;
33438: pixelout<=1'b1;
33439: pixelout<=1'b1;
33440: pixelout<=1'b1;
33441: pixelout<=1'b1;
33442: pixelout<=1'b1;
33443: pixelout<=1'b1;
33444: pixelout<=1'b1;
33445: pixelout<=1'b1;
33446: pixelout<=1'b1;
33447: pixelout<=1'b1;
33448: pixelout<=1'b1;
33449: pixelout<=1'b1;
33450: pixelout<=1'b1;
33451: pixelout<=1'b1;
33452: pixelout<=1'b1;
33453: pixelout<=1'b1;
33454: pixelout<=1'b1;
33455: pixelout<=1'b1;
33456: pixelout<=1'b1;
33457: pixelout<=1'b1;
33458: pixelout<=1'b1;
33459: pixelout<=1'b1;
33460: pixelout<=1'b1;
33461: pixelout<=1'b1;
33462: pixelout<=1'b1;
33463: pixelout<=1'b1;
33464: pixelout<=1'b1;
33465: pixelout<=1'b1;
33466: pixelout<=1'b1;
33467: pixelout<=1'b1;
33468: pixelout<=1'b1;
33469: pixelout<=1'b1;
33470: pixelout<=1'b1;
33471: pixelout<=1'b1;
33472: pixelout<=1'b1;
33473: pixelout<=1'b1;
33474: pixelout<=1'b1;
33475: pixelout<=1'b1;
33476: pixelout<=1'b1;
33477: pixelout<=1'b1;
33478: pixelout<=1'b1;
33479: pixelout<=1'b1;
33480: pixelout<=1'b1;
33481: pixelout<=1'b1;
33482: pixelout<=1'b1;
33483: pixelout<=1'b1;
33484: pixelout<=1'b1;
33485: pixelout<=1'b1;
33486: pixelout<=1'b1;
33487: pixelout<=1'b1;
33488: pixelout<=1'b1;
33489: pixelout<=1'b1;
33490: pixelout<=1'b1;
33491: pixelout<=1'b1;
33492: pixelout<=1'b1;
33493: pixelout<=1'b1;
33494: pixelout<=1'b1;
33495: pixelout<=1'b1;
33496: pixelout<=1'b1;
33497: pixelout<=1'b1;
33498: pixelout<=1'b1;
33499: pixelout<=1'b1;
33500: pixelout<=1'b1;
33501: pixelout<=1'b1;
33502: pixelout<=1'b1;
33503: pixelout<=1'b1;
33504: pixelout<=1'b1;
33505: pixelout<=1'b1;
33506: pixelout<=1'b1;
33507: pixelout<=1'b0;
33508: pixelout<=1'b0;
33509: pixelout<=1'b0;
33510: pixelout<=1'b0;
33511: pixelout<=1'b1;
33512: pixelout<=1'b1;
33513: pixelout<=1'b1;
33514: pixelout<=1'b1;
33515: pixelout<=1'b1;
33516: pixelout<=1'b1;
33517: pixelout<=1'b1;
33518: pixelout<=1'b1;
33519: pixelout<=1'b1;
33520: pixelout<=1'b1;
33521: pixelout<=1'b1;
33522: pixelout<=1'b1;
33523: pixelout<=1'b1;
33524: pixelout<=1'b1;
33525: pixelout<=1'b1;
33526: pixelout<=1'b1;
33527: pixelout<=1'b1;
33528: pixelout<=1'b1;
33529: pixelout<=1'b1;
33530: pixelout<=1'b1;
33531: pixelout<=1'b1;
33532: pixelout<=1'b1;
33533: pixelout<=1'b1;
33534: pixelout<=1'b1;
33535: pixelout<=1'b1;
33536: pixelout<=1'b1;
33537: pixelout<=1'b1;
33538: pixelout<=1'b1;
33539: pixelout<=1'b1;
33540: pixelout<=1'b1;
33541: pixelout<=1'b1;
33542: pixelout<=1'b1;
33543: pixelout<=1'b1;
33544: pixelout<=1'b1;
33545: pixelout<=1'b1;
33546: pixelout<=1'b1;
33547: pixelout<=1'b1;
33548: pixelout<=1'b1;
33549: pixelout<=1'b1;
33550: pixelout<=1'b1;
33551: pixelout<=1'b1;
33552: pixelout<=1'b1;
33553: pixelout<=1'b0;
33554: pixelout<=1'b0;
33555: pixelout<=1'b0;
33556: pixelout<=1'b0;
33557: pixelout<=1'b1;
33558: pixelout<=1'b1;
33559: pixelout<=1'b1;
33560: pixelout<=1'b1;
33561: pixelout<=1'b1;
33562: pixelout<=1'b1;
33563: pixelout<=1'b1;
33564: pixelout<=1'b1;
33565: pixelout<=1'b1;
33566: pixelout<=1'b1;
33567: pixelout<=1'b1;
33568: pixelout<=1'b1;
33569: pixelout<=1'b1;
33570: pixelout<=1'b1;
33571: pixelout<=1'b1;
33572: pixelout<=1'b1;
33573: pixelout<=1'b1;
33574: pixelout<=1'b1;
33575: pixelout<=1'b1;
33576: pixelout<=1'b1;
33577: pixelout<=1'b1;
33578: pixelout<=1'b1;
33579: pixelout<=1'b1;
33580: pixelout<=1'b1;
33581: pixelout<=1'b1;
33582: pixelout<=1'b1;
33583: pixelout<=1'b1;
33584: pixelout<=1'b1;
33585: pixelout<=1'b1;
33586: pixelout<=1'b1;
33587: pixelout<=1'b1;
33588: pixelout<=1'b1;
33589: pixelout<=1'b1;
33590: pixelout<=1'b1;
33591: pixelout<=1'b1;
33592: pixelout<=1'b1;
33593: pixelout<=1'b1;
33594: pixelout<=1'b1;
33595: pixelout<=1'b1;
33596: pixelout<=1'b1;
33597: pixelout<=1'b1;
33598: pixelout<=1'b1;
33599: pixelout<=1'b1;
33600: pixelout<=1'b1;
33601: pixelout<=1'b1;
33602: pixelout<=1'b1;
33603: pixelout<=1'b1;
33604: pixelout<=1'b1;
33605: pixelout<=1'b1;
33606: pixelout<=1'b1;
33607: pixelout<=1'b1;
33608: pixelout<=1'b1;
33609: pixelout<=1'b1;
33610: pixelout<=1'b1;
33611: pixelout<=1'b1;
33612: pixelout<=1'b1;
33613: pixelout<=1'b1;
33614: pixelout<=1'b1;
33615: pixelout<=1'b1;
33616: pixelout<=1'b1;
33617: pixelout<=1'b1;
33618: pixelout<=1'b1;
33619: pixelout<=1'b1;
33620: pixelout<=1'b1;
33621: pixelout<=1'b1;
33622: pixelout<=1'b1;
33623: pixelout<=1'b1;
33624: pixelout<=1'b1;
33625: pixelout<=1'b1;
33626: pixelout<=1'b1;
33627: pixelout<=1'b1;
33628: pixelout<=1'b1;
33629: pixelout<=1'b1;
33630: pixelout<=1'b1;
33631: pixelout<=1'b1;
33632: pixelout<=1'b1;
33633: pixelout<=1'b1;
33634: pixelout<=1'b1;
33635: pixelout<=1'b1;
33636: pixelout<=1'b1;
33637: pixelout<=1'b1;
33638: pixelout<=1'b1;
33639: pixelout<=1'b1;
33640: pixelout<=1'b1;
33641: pixelout<=1'b1;
33642: pixelout<=1'b1;
33643: pixelout<=1'b1;
33644: pixelout<=1'b1;
33645: pixelout<=1'b1;
33646: pixelout<=1'b1;
33647: pixelout<=1'b1;
33648: pixelout<=1'b1;
33649: pixelout<=1'b1;
33650: pixelout<=1'b1;
33651: pixelout<=1'b1;
33652: pixelout<=1'b1;
33653: pixelout<=1'b1;
33654: pixelout<=1'b1;
33655: pixelout<=1'b1;
33656: pixelout<=1'b1;
33657: pixelout<=1'b1;
33658: pixelout<=1'b1;
33659: pixelout<=1'b1;
33660: pixelout<=1'b1;
33661: pixelout<=1'b1;
33662: pixelout<=1'b1;
33663: pixelout<=1'b1;
33664: pixelout<=1'b1;
33665: pixelout<=1'b1;
33666: pixelout<=1'b1;
33667: pixelout<=1'b1;
33668: pixelout<=1'b1;
33669: pixelout<=1'b1;
33670: pixelout<=1'b1;
33671: pixelout<=1'b1;
33672: pixelout<=1'b1;
33673: pixelout<=1'b1;
33674: pixelout<=1'b1;
33675: pixelout<=1'b1;
33676: pixelout<=1'b1;
33677: pixelout<=1'b1;
33678: pixelout<=1'b1;
33679: pixelout<=1'b1;
33680: pixelout<=1'b1;
33681: pixelout<=1'b1;
33682: pixelout<=1'b1;
33683: pixelout<=1'b1;
33684: pixelout<=1'b1;
33685: pixelout<=1'b1;
33686: pixelout<=1'b1;
33687: pixelout<=1'b1;
33688: pixelout<=1'b1;
33689: pixelout<=1'b1;
33690: pixelout<=1'b1;
33691: pixelout<=1'b1;
33692: pixelout<=1'b1;
33693: pixelout<=1'b1;
33694: pixelout<=1'b1;
33695: pixelout<=1'b1;
33696: pixelout<=1'b1;
33697: pixelout<=1'b1;
33698: pixelout<=1'b1;
33699: pixelout<=1'b1;
33700: pixelout<=1'b1;
33701: pixelout<=1'b1;
33702: pixelout<=1'b1;
33703: pixelout<=1'b1;
33704: pixelout<=1'b1;
33705: pixelout<=1'b1;
33706: pixelout<=1'b1;
33707: pixelout<=1'b1;
33708: pixelout<=1'b1;
33709: pixelout<=1'b1;
33710: pixelout<=1'b1;
33711: pixelout<=1'b1;
33712: pixelout<=1'b1;
33713: pixelout<=1'b1;
33714: pixelout<=1'b1;
33715: pixelout<=1'b1;
33716: pixelout<=1'b1;
33717: pixelout<=1'b1;
33718: pixelout<=1'b1;
33719: pixelout<=1'b1;
33720: pixelout<=1'b1;
33721: pixelout<=1'b1;
33722: pixelout<=1'b1;
33723: pixelout<=1'b1;
33724: pixelout<=1'b1;
33725: pixelout<=1'b1;
33726: pixelout<=1'b1;
33727: pixelout<=1'b1;
33728: pixelout<=1'b1;
33729: pixelout<=1'b1;
33730: pixelout<=1'b1;
33731: pixelout<=1'b1;
33732: pixelout<=1'b1;
33733: pixelout<=1'b1;
33734: pixelout<=1'b1;
33735: pixelout<=1'b1;
33736: pixelout<=1'b1;
33737: pixelout<=1'b1;
33738: pixelout<=1'b1;
33739: pixelout<=1'b1;
33740: pixelout<=1'b1;
33741: pixelout<=1'b1;
33742: pixelout<=1'b1;
33743: pixelout<=1'b1;
33744: pixelout<=1'b1;
33745: pixelout<=1'b1;
33746: pixelout<=1'b1;
33747: pixelout<=1'b1;
33748: pixelout<=1'b1;
33749: pixelout<=1'b1;
33750: pixelout<=1'b1;
33751: pixelout<=1'b1;
33752: pixelout<=1'b1;
33753: pixelout<=1'b1;
33754: pixelout<=1'b1;
33755: pixelout<=1'b1;
33756: pixelout<=1'b1;
33757: pixelout<=1'b1;
33758: pixelout<=1'b1;
33759: pixelout<=1'b1;
33760: pixelout<=1'b1;
33761: pixelout<=1'b1;
33762: pixelout<=1'b1;
33763: pixelout<=1'b1;
33764: pixelout<=1'b1;
33765: pixelout<=1'b1;
33766: pixelout<=1'b1;
33767: pixelout<=1'b1;
33768: pixelout<=1'b1;
33769: pixelout<=1'b1;
33770: pixelout<=1'b1;
33771: pixelout<=1'b1;
33772: pixelout<=1'b1;
33773: pixelout<=1'b1;
33774: pixelout<=1'b1;
33775: pixelout<=1'b1;
33776: pixelout<=1'b1;
33777: pixelout<=1'b1;
33778: pixelout<=1'b1;
33779: pixelout<=1'b1;
33780: pixelout<=1'b1;
33781: pixelout<=1'b1;
33782: pixelout<=1'b1;
33783: pixelout<=1'b1;
33784: pixelout<=1'b1;
33785: pixelout<=1'b1;
33786: pixelout<=1'b1;
33787: pixelout<=1'b1;
33788: pixelout<=1'b1;
33789: pixelout<=1'b1;
33790: pixelout<=1'b1;
33791: pixelout<=1'b1;
33792: pixelout<=1'b1;
33793: pixelout<=1'b1;
33794: pixelout<=1'b1;
33795: pixelout<=1'b1;
33796: pixelout<=1'b1;
33797: pixelout<=1'b1;
33798: pixelout<=1'b1;
33799: pixelout<=1'b1;
33800: pixelout<=1'b1;
33801: pixelout<=1'b1;
33802: pixelout<=1'b1;
33803: pixelout<=1'b1;
33804: pixelout<=1'b1;
33805: pixelout<=1'b1;
33806: pixelout<=1'b1;
33807: pixelout<=1'b1;
33808: pixelout<=1'b1;
33809: pixelout<=1'b1;
33810: pixelout<=1'b1;
33811: pixelout<=1'b1;
33812: pixelout<=1'b1;
33813: pixelout<=1'b1;
33814: pixelout<=1'b1;
33815: pixelout<=1'b1;
33816: pixelout<=1'b1;
33817: pixelout<=1'b1;
33818: pixelout<=1'b1;
33819: pixelout<=1'b1;
33820: pixelout<=1'b1;
33821: pixelout<=1'b1;
33822: pixelout<=1'b1;
33823: pixelout<=1'b1;
33824: pixelout<=1'b1;
33825: pixelout<=1'b1;
33826: pixelout<=1'b1;
33827: pixelout<=1'b1;
33828: pixelout<=1'b1;
33829: pixelout<=1'b1;
33830: pixelout<=1'b1;
33831: pixelout<=1'b1;
33832: pixelout<=1'b1;
33833: pixelout<=1'b1;
33834: pixelout<=1'b1;
33835: pixelout<=1'b1;
33836: pixelout<=1'b1;
33837: pixelout<=1'b1;
33838: pixelout<=1'b1;
33839: pixelout<=1'b1;
33840: pixelout<=1'b1;
33841: pixelout<=1'b1;
33842: pixelout<=1'b1;
33843: pixelout<=1'b1;
33844: pixelout<=1'b1;
33845: pixelout<=1'b1;
33846: pixelout<=1'b1;
33847: pixelout<=1'b1;
33848: pixelout<=1'b1;
33849: pixelout<=1'b1;
33850: pixelout<=1'b1;
33851: pixelout<=1'b1;
33852: pixelout<=1'b1;
33853: pixelout<=1'b1;
33854: pixelout<=1'b1;
33855: pixelout<=1'b1;
33856: pixelout<=1'b1;
33857: pixelout<=1'b1;
33858: pixelout<=1'b1;
33859: pixelout<=1'b1;
33860: pixelout<=1'b1;
33861: pixelout<=1'b1;
33862: pixelout<=1'b1;
33863: pixelout<=1'b1;
33864: pixelout<=1'b1;
33865: pixelout<=1'b1;
33866: pixelout<=1'b1;
33867: pixelout<=1'b1;
33868: pixelout<=1'b1;
33869: pixelout<=1'b1;
33870: pixelout<=1'b1;
33871: pixelout<=1'b1;
33872: pixelout<=1'b1;
33873: pixelout<=1'b1;
33874: pixelout<=1'b1;
33875: pixelout<=1'b1;
33876: pixelout<=1'b1;
33877: pixelout<=1'b1;
33878: pixelout<=1'b1;
33879: pixelout<=1'b1;
33880: pixelout<=1'b1;
33881: pixelout<=1'b1;
33882: pixelout<=1'b1;
33883: pixelout<=1'b1;
33884: pixelout<=1'b1;
33885: pixelout<=1'b1;
33886: pixelout<=1'b1;
33887: pixelout<=1'b1;
33888: pixelout<=1'b1;
33889: pixelout<=1'b1;
33890: pixelout<=1'b1;
33891: pixelout<=1'b1;
33892: pixelout<=1'b1;
33893: pixelout<=1'b1;
33894: pixelout<=1'b1;
33895: pixelout<=1'b1;
33896: pixelout<=1'b1;
33897: pixelout<=1'b1;
33898: pixelout<=1'b1;
33899: pixelout<=1'b1;
33900: pixelout<=1'b1;
33901: pixelout<=1'b1;
33902: pixelout<=1'b1;
33903: pixelout<=1'b1;
33904: pixelout<=1'b1;
33905: pixelout<=1'b1;
33906: pixelout<=1'b1;
33907: pixelout<=1'b1;
33908: pixelout<=1'b1;
33909: pixelout<=1'b1;
33910: pixelout<=1'b1;
33911: pixelout<=1'b1;
33912: pixelout<=1'b1;
33913: pixelout<=1'b1;
33914: pixelout<=1'b1;
33915: pixelout<=1'b1;
33916: pixelout<=1'b1;
33917: pixelout<=1'b1;
33918: pixelout<=1'b1;
33919: pixelout<=1'b1;
33920: pixelout<=1'b1;
33921: pixelout<=1'b1;
33922: pixelout<=1'b1;
33923: pixelout<=1'b1;
33924: pixelout<=1'b1;
33925: pixelout<=1'b1;
33926: pixelout<=1'b1;
33927: pixelout<=1'b1;
33928: pixelout<=1'b1;
33929: pixelout<=1'b1;
33930: pixelout<=1'b1;
33931: pixelout<=1'b1;
33932: pixelout<=1'b1;
33933: pixelout<=1'b1;
33934: pixelout<=1'b1;
33935: pixelout<=1'b1;
33936: pixelout<=1'b1;
33937: pixelout<=1'b1;
33938: pixelout<=1'b1;
33939: pixelout<=1'b1;
33940: pixelout<=1'b1;
33941: pixelout<=1'b1;
33942: pixelout<=1'b1;
33943: pixelout<=1'b1;
33944: pixelout<=1'b1;
33945: pixelout<=1'b1;
33946: pixelout<=1'b1;
33947: pixelout<=1'b1;
33948: pixelout<=1'b1;
33949: pixelout<=1'b1;
33950: pixelout<=1'b1;
33951: pixelout<=1'b1;
33952: pixelout<=1'b1;
33953: pixelout<=1'b1;
33954: pixelout<=1'b1;
33955: pixelout<=1'b1;
33956: pixelout<=1'b1;
33957: pixelout<=1'b1;
33958: pixelout<=1'b1;
33959: pixelout<=1'b1;
33960: pixelout<=1'b1;
33961: pixelout<=1'b1;
33962: pixelout<=1'b1;
33963: pixelout<=1'b1;
33964: pixelout<=1'b1;
33965: pixelout<=1'b1;
33966: pixelout<=1'b1;
33967: pixelout<=1'b1;
33968: pixelout<=1'b1;
33969: pixelout<=1'b1;
33970: pixelout<=1'b1;
33971: pixelout<=1'b1;
33972: pixelout<=1'b1;
33973: pixelout<=1'b1;
33974: pixelout<=1'b1;
33975: pixelout<=1'b1;
33976: pixelout<=1'b1;
33977: pixelout<=1'b1;
33978: pixelout<=1'b1;
33979: pixelout<=1'b1;
33980: pixelout<=1'b1;
33981: pixelout<=1'b1;
33982: pixelout<=1'b1;
33983: pixelout<=1'b1;
33984: pixelout<=1'b1;
33985: pixelout<=1'b1;
33986: pixelout<=1'b1;
33987: pixelout<=1'b1;
33988: pixelout<=1'b1;
33989: pixelout<=1'b1;
33990: pixelout<=1'b1;
33991: pixelout<=1'b1;
33992: pixelout<=1'b1;
33993: pixelout<=1'b1;
33994: pixelout<=1'b1;
33995: pixelout<=1'b1;
33996: pixelout<=1'b1;
33997: pixelout<=1'b1;
33998: pixelout<=1'b1;
33999: pixelout<=1'b1;
34000: pixelout<=1'b1;
34001: pixelout<=1'b1;
34002: pixelout<=1'b1;
34003: pixelout<=1'b1;
34004: pixelout<=1'b1;
34005: pixelout<=1'b1;
34006: pixelout<=1'b1;
34007: pixelout<=1'b1;
34008: pixelout<=1'b1;
34009: pixelout<=1'b1;
34010: pixelout<=1'b1;
34011: pixelout<=1'b1;
34012: pixelout<=1'b1;
34013: pixelout<=1'b1;
34014: pixelout<=1'b1;
34015: pixelout<=1'b1;
34016: pixelout<=1'b1;
34017: pixelout<=1'b1;
34018: pixelout<=1'b1;
34019: pixelout<=1'b1;
34020: pixelout<=1'b1;
34021: pixelout<=1'b1;
34022: pixelout<=1'b1;
34023: pixelout<=1'b1;
34024: pixelout<=1'b1;
34025: pixelout<=1'b1;
34026: pixelout<=1'b1;
34027: pixelout<=1'b1;
34028: pixelout<=1'b1;
34029: pixelout<=1'b1;
34030: pixelout<=1'b1;
34031: pixelout<=1'b1;
34032: pixelout<=1'b1;
34033: pixelout<=1'b1;
34034: pixelout<=1'b1;
34035: pixelout<=1'b1;
34036: pixelout<=1'b1;
34037: pixelout<=1'b1;
34038: pixelout<=1'b1;
34039: pixelout<=1'b1;
34040: pixelout<=1'b1;
34041: pixelout<=1'b1;
34042: pixelout<=1'b1;
34043: pixelout<=1'b1;
34044: pixelout<=1'b1;
34045: pixelout<=1'b1;
34046: pixelout<=1'b1;
34047: pixelout<=1'b1;
34048: pixelout<=1'b1;
34049: pixelout<=1'b1;
34050: pixelout<=1'b1;
34051: pixelout<=1'b1;
34052: pixelout<=1'b1;
34053: pixelout<=1'b1;
34054: pixelout<=1'b1;
34055: pixelout<=1'b1;
34056: pixelout<=1'b1;
34057: pixelout<=1'b1;
34058: pixelout<=1'b1;
34059: pixelout<=1'b1;
34060: pixelout<=1'b1;
34061: pixelout<=1'b1;
34062: pixelout<=1'b1;
34063: pixelout<=1'b1;
34064: pixelout<=1'b1;
34065: pixelout<=1'b1;
34066: pixelout<=1'b1;
34067: pixelout<=1'b1;
34068: pixelout<=1'b1;
34069: pixelout<=1'b1;
34070: pixelout<=1'b1;
34071: pixelout<=1'b1;
34072: pixelout<=1'b1;
34073: pixelout<=1'b1;
34074: pixelout<=1'b1;
34075: pixelout<=1'b1;
34076: pixelout<=1'b1;
34077: pixelout<=1'b1;
34078: pixelout<=1'b1;
34079: pixelout<=1'b1;
34080: pixelout<=1'b1;
34081: pixelout<=1'b1;
34082: pixelout<=1'b1;
34083: pixelout<=1'b1;
34084: pixelout<=1'b1;
34085: pixelout<=1'b1;
34086: pixelout<=1'b1;
34087: pixelout<=1'b1;
34088: pixelout<=1'b1;
34089: pixelout<=1'b1;
34090: pixelout<=1'b1;
34091: pixelout<=1'b1;
34092: pixelout<=1'b1;
34093: pixelout<=1'b1;
34094: pixelout<=1'b1;
34095: pixelout<=1'b1;
34096: pixelout<=1'b1;
34097: pixelout<=1'b1;
34098: pixelout<=1'b1;
34099: pixelout<=1'b1;
34100: pixelout<=1'b1;
34101: pixelout<=1'b1;
34102: pixelout<=1'b1;
34103: pixelout<=1'b1;
34104: pixelout<=1'b1;
34105: pixelout<=1'b1;
34106: pixelout<=1'b1;
34107: pixelout<=1'b1;
34108: pixelout<=1'b1;
34109: pixelout<=1'b1;
34110: pixelout<=1'b1;
34111: pixelout<=1'b1;
34112: pixelout<=1'b1;
34113: pixelout<=1'b1;
34114: pixelout<=1'b1;
34115: pixelout<=1'b1;
34116: pixelout<=1'b1;
34117: pixelout<=1'b1;
34118: pixelout<=1'b1;
34119: pixelout<=1'b1;
34120: pixelout<=1'b1;
34121: pixelout<=1'b1;
34122: pixelout<=1'b1;
34123: pixelout<=1'b1;
34124: pixelout<=1'b1;
34125: pixelout<=1'b1;
34126: pixelout<=1'b1;
34127: pixelout<=1'b1;
34128: pixelout<=1'b1;
34129: pixelout<=1'b1;
34130: pixelout<=1'b1;
34131: pixelout<=1'b1;
34132: pixelout<=1'b1;
34133: pixelout<=1'b1;
34134: pixelout<=1'b1;
34135: pixelout<=1'b1;
34136: pixelout<=1'b1;
34137: pixelout<=1'b1;
34138: pixelout<=1'b1;
34139: pixelout<=1'b1;
34140: pixelout<=1'b1;
34141: pixelout<=1'b1;
34142: pixelout<=1'b1;
34143: pixelout<=1'b1;
34144: pixelout<=1'b1;
34145: pixelout<=1'b1;
34146: pixelout<=1'b1;
34147: pixelout<=1'b1;
34148: pixelout<=1'b1;
34149: pixelout<=1'b1;
34150: pixelout<=1'b1;
34151: pixelout<=1'b1;
34152: pixelout<=1'b1;
34153: pixelout<=1'b1;
34154: pixelout<=1'b1;
34155: pixelout<=1'b1;
34156: pixelout<=1'b1;
34157: pixelout<=1'b1;
34158: pixelout<=1'b1;
34159: pixelout<=1'b1;
34160: pixelout<=1'b1;
34161: pixelout<=1'b1;
34162: pixelout<=1'b1;
34163: pixelout<=1'b1;
34164: pixelout<=1'b1;
34165: pixelout<=1'b1;
34166: pixelout<=1'b1;
34167: pixelout<=1'b1;
34168: pixelout<=1'b1;
34169: pixelout<=1'b1;
34170: pixelout<=1'b1;
34171: pixelout<=1'b1;
34172: pixelout<=1'b1;
34173: pixelout<=1'b1;
34174: pixelout<=1'b1;
34175: pixelout<=1'b1;
34176: pixelout<=1'b1;
34177: pixelout<=1'b1;
34178: pixelout<=1'b1;
34179: pixelout<=1'b1;
34180: pixelout<=1'b1;
34181: pixelout<=1'b1;
34182: pixelout<=1'b1;
34183: pixelout<=1'b1;
34184: pixelout<=1'b1;
34185: pixelout<=1'b1;
34186: pixelout<=1'b1;
34187: pixelout<=1'b1;
34188: pixelout<=1'b1;
34189: pixelout<=1'b1;
34190: pixelout<=1'b1;
34191: pixelout<=1'b1;
34192: pixelout<=1'b1;
34193: pixelout<=1'b1;
34194: pixelout<=1'b1;
34195: pixelout<=1'b1;
34196: pixelout<=1'b1;
34197: pixelout<=1'b1;
34198: pixelout<=1'b1;
34199: pixelout<=1'b1;
34200: pixelout<=1'b1;
34201: pixelout<=1'b1;
34202: pixelout<=1'b1;
34203: pixelout<=1'b1;
34204: pixelout<=1'b1;
34205: pixelout<=1'b1;
34206: pixelout<=1'b1;
34207: pixelout<=1'b1;
34208: pixelout<=1'b1;
34209: pixelout<=1'b1;
34210: pixelout<=1'b1;
34211: pixelout<=1'b1;
34212: pixelout<=1'b1;
34213: pixelout<=1'b1;
34214: pixelout<=1'b1;
34215: pixelout<=1'b1;
34216: pixelout<=1'b1;
34217: pixelout<=1'b1;
34218: pixelout<=1'b1;
34219: pixelout<=1'b1;
34220: pixelout<=1'b1;
34221: pixelout<=1'b1;
34222: pixelout<=1'b1;
34223: pixelout<=1'b1;
34224: pixelout<=1'b1;
34225: pixelout<=1'b1;
34226: pixelout<=1'b1;
34227: pixelout<=1'b1;
34228: pixelout<=1'b1;
34229: pixelout<=1'b1;
34230: pixelout<=1'b1;
34231: pixelout<=1'b1;
34232: pixelout<=1'b1;
34233: pixelout<=1'b1;
34234: pixelout<=1'b1;
34235: pixelout<=1'b1;
34236: pixelout<=1'b1;
34237: pixelout<=1'b1;
34238: pixelout<=1'b1;
34239: pixelout<=1'b1;
34240: pixelout<=1'b1;
34241: pixelout<=1'b1;
34242: pixelout<=1'b1;
34243: pixelout<=1'b1;
34244: pixelout<=1'b1;
34245: pixelout<=1'b1;
34246: pixelout<=1'b1;
34247: pixelout<=1'b1;
34248: pixelout<=1'b1;
34249: pixelout<=1'b1;
34250: pixelout<=1'b1;
34251: pixelout<=1'b1;
34252: pixelout<=1'b1;
34253: pixelout<=1'b1;
34254: pixelout<=1'b1;
34255: pixelout<=1'b1;
34256: pixelout<=1'b1;
34257: pixelout<=1'b1;
34258: pixelout<=1'b1;
34259: pixelout<=1'b1;
34260: pixelout<=1'b1;
34261: pixelout<=1'b1;
34262: pixelout<=1'b1;
34263: pixelout<=1'b1;
34264: pixelout<=1'b1;
34265: pixelout<=1'b1;
34266: pixelout<=1'b1;
34267: pixelout<=1'b1;
34268: pixelout<=1'b1;
34269: pixelout<=1'b1;
34270: pixelout<=1'b1;
34271: pixelout<=1'b1;
34272: pixelout<=1'b1;
34273: pixelout<=1'b1;
34274: pixelout<=1'b1;
34275: pixelout<=1'b1;
34276: pixelout<=1'b1;
34277: pixelout<=1'b1;
34278: pixelout<=1'b1;
34279: pixelout<=1'b1;
34280: pixelout<=1'b1;
34281: pixelout<=1'b1;
34282: pixelout<=1'b1;
34283: pixelout<=1'b1;
34284: pixelout<=1'b1;
34285: pixelout<=1'b1;
34286: pixelout<=1'b1;
34287: pixelout<=1'b1;
34288: pixelout<=1'b1;
34289: pixelout<=1'b1;
34290: pixelout<=1'b1;
34291: pixelout<=1'b1;
34292: pixelout<=1'b1;
34293: pixelout<=1'b1;
34294: pixelout<=1'b1;
34295: pixelout<=1'b1;
34296: pixelout<=1'b1;
34297: pixelout<=1'b1;
34298: pixelout<=1'b1;
34299: pixelout<=1'b1;
34300: pixelout<=1'b1;
34301: pixelout<=1'b1;
34302: pixelout<=1'b1;
34303: pixelout<=1'b1;
34304: pixelout<=1'b1;
34305: pixelout<=1'b1;
34306: pixelout<=1'b1;
34307: pixelout<=1'b1;
34308: pixelout<=1'b1;
34309: pixelout<=1'b1;
34310: pixelout<=1'b1;
34311: pixelout<=1'b1;
34312: pixelout<=1'b1;
34313: pixelout<=1'b1;
34314: pixelout<=1'b1;
34315: pixelout<=1'b1;
34316: pixelout<=1'b1;
34317: pixelout<=1'b1;
34318: pixelout<=1'b1;
34319: pixelout<=1'b1;
34320: pixelout<=1'b1;
34321: pixelout<=1'b1;
34322: pixelout<=1'b1;
34323: pixelout<=1'b1;
34324: pixelout<=1'b1;
34325: pixelout<=1'b1;
34326: pixelout<=1'b1;
34327: pixelout<=1'b1;
34328: pixelout<=1'b1;
34329: pixelout<=1'b1;
34330: pixelout<=1'b1;
34331: pixelout<=1'b1;
34332: pixelout<=1'b1;
34333: pixelout<=1'b1;
34334: pixelout<=1'b1;
34335: pixelout<=1'b1;
34336: pixelout<=1'b1;
34337: pixelout<=1'b1;
34338: pixelout<=1'b1;
34339: pixelout<=1'b1;
34340: pixelout<=1'b1;
34341: pixelout<=1'b1;
34342: pixelout<=1'b1;
34343: pixelout<=1'b1;
34344: pixelout<=1'b1;
34345: pixelout<=1'b1;
34346: pixelout<=1'b1;
34347: pixelout<=1'b1;
34348: pixelout<=1'b1;
34349: pixelout<=1'b1;
34350: pixelout<=1'b1;
34351: pixelout<=1'b1;
34352: pixelout<=1'b1;
34353: pixelout<=1'b1;
34354: pixelout<=1'b1;
34355: pixelout<=1'b1;
34356: pixelout<=1'b1;
34357: pixelout<=1'b1;
34358: pixelout<=1'b1;
34359: pixelout<=1'b1;
34360: pixelout<=1'b1;
34361: pixelout<=1'b1;
34362: pixelout<=1'b1;
34363: pixelout<=1'b1;
34364: pixelout<=1'b1;
34365: pixelout<=1'b1;
34366: pixelout<=1'b1;
34367: pixelout<=1'b1;
34368: pixelout<=1'b1;
34369: pixelout<=1'b1;
34370: pixelout<=1'b1;
34371: pixelout<=1'b1;
34372: pixelout<=1'b1;
34373: pixelout<=1'b1;
34374: pixelout<=1'b1;
34375: pixelout<=1'b1;
34376: pixelout<=1'b1;
34377: pixelout<=1'b1;
34378: pixelout<=1'b1;
34379: pixelout<=1'b1;
34380: pixelout<=1'b1;
34381: pixelout<=1'b1;
34382: pixelout<=1'b1;
34383: pixelout<=1'b1;
34384: pixelout<=1'b1;
34385: pixelout<=1'b1;
34386: pixelout<=1'b1;
34387: pixelout<=1'b1;
34388: pixelout<=1'b1;
34389: pixelout<=1'b1;
34390: pixelout<=1'b1;
34391: pixelout<=1'b1;
34392: pixelout<=1'b1;
34393: pixelout<=1'b1;
34394: pixelout<=1'b1;
34395: pixelout<=1'b1;
34396: pixelout<=1'b1;
34397: pixelout<=1'b1;
34398: pixelout<=1'b1;
34399: pixelout<=1'b1;
34400: pixelout<=1'b1;
34401: pixelout<=1'b1;
34402: pixelout<=1'b1;
34403: pixelout<=1'b1;
34404: pixelout<=1'b1;
34405: pixelout<=1'b1;
34406: pixelout<=1'b1;
34407: pixelout<=1'b1;
34408: pixelout<=1'b1;
34409: pixelout<=1'b1;
34410: pixelout<=1'b1;
34411: pixelout<=1'b1;
34412: pixelout<=1'b1;
34413: pixelout<=1'b1;
34414: pixelout<=1'b1;
34415: pixelout<=1'b1;
34416: pixelout<=1'b1;
34417: pixelout<=1'b1;
34418: pixelout<=1'b1;
34419: pixelout<=1'b1;
34420: pixelout<=1'b1;
34421: pixelout<=1'b1;
34422: pixelout<=1'b1;
34423: pixelout<=1'b1;
34424: pixelout<=1'b1;
34425: pixelout<=1'b1;
34426: pixelout<=1'b1;
34427: pixelout<=1'b1;
34428: pixelout<=1'b1;
34429: pixelout<=1'b1;
34430: pixelout<=1'b1;
34431: pixelout<=1'b1;
34432: pixelout<=1'b1;
34433: pixelout<=1'b1;
34434: pixelout<=1'b1;
34435: pixelout<=1'b1;
34436: pixelout<=1'b1;
34437: pixelout<=1'b1;
34438: pixelout<=1'b1;
34439: pixelout<=1'b1;
34440: pixelout<=1'b1;
34441: pixelout<=1'b1;
34442: pixelout<=1'b1;
34443: pixelout<=1'b1;
34444: pixelout<=1'b1;
34445: pixelout<=1'b1;
34446: pixelout<=1'b1;
34447: pixelout<=1'b1;
34448: pixelout<=1'b1;
34449: pixelout<=1'b1;
34450: pixelout<=1'b1;
34451: pixelout<=1'b1;
34452: pixelout<=1'b1;
34453: pixelout<=1'b1;
34454: pixelout<=1'b1;
34455: pixelout<=1'b1;
34456: pixelout<=1'b1;
34457: pixelout<=1'b1;
34458: pixelout<=1'b1;
34459: pixelout<=1'b1;
34460: pixelout<=1'b1;
34461: pixelout<=1'b1;
34462: pixelout<=1'b1;
34463: pixelout<=1'b1;
34464: pixelout<=1'b1;
34465: pixelout<=1'b1;
34466: pixelout<=1'b1;
34467: pixelout<=1'b1;
34468: pixelout<=1'b1;
34469: pixelout<=1'b1;
34470: pixelout<=1'b1;
34471: pixelout<=1'b1;
34472: pixelout<=1'b1;
34473: pixelout<=1'b1;
34474: pixelout<=1'b1;
34475: pixelout<=1'b1;
34476: pixelout<=1'b1;
34477: pixelout<=1'b1;
34478: pixelout<=1'b1;
34479: pixelout<=1'b1;
34480: pixelout<=1'b1;
34481: pixelout<=1'b1;
34482: pixelout<=1'b1;
34483: pixelout<=1'b1;
34484: pixelout<=1'b1;
34485: pixelout<=1'b1;
34486: pixelout<=1'b1;
34487: pixelout<=1'b1;
34488: pixelout<=1'b1;
34489: pixelout<=1'b1;
34490: pixelout<=1'b1;
34491: pixelout<=1'b1;
34492: pixelout<=1'b1;
34493: pixelout<=1'b1;
34494: pixelout<=1'b1;
34495: pixelout<=1'b1;
34496: pixelout<=1'b1;
34497: pixelout<=1'b1;
34498: pixelout<=1'b1;
34499: pixelout<=1'b1;
34500: pixelout<=1'b1;
34501: pixelout<=1'b1;
34502: pixelout<=1'b1;
34503: pixelout<=1'b1;
34504: pixelout<=1'b1;
34505: pixelout<=1'b1;
34506: pixelout<=1'b1;
34507: pixelout<=1'b1;
34508: pixelout<=1'b1;
34509: pixelout<=1'b1;
34510: pixelout<=1'b1;
34511: pixelout<=1'b1;
34512: pixelout<=1'b1;
34513: pixelout<=1'b1;
34514: pixelout<=1'b1;
34515: pixelout<=1'b1;
34516: pixelout<=1'b1;
34517: pixelout<=1'b1;
34518: pixelout<=1'b1;
34519: pixelout<=1'b1;
34520: pixelout<=1'b1;
34521: pixelout<=1'b1;
34522: pixelout<=1'b1;
34523: pixelout<=1'b1;
34524: pixelout<=1'b1;
34525: pixelout<=1'b1;
34526: pixelout<=1'b1;
34527: pixelout<=1'b1;
34528: pixelout<=1'b1;
34529: pixelout<=1'b1;
34530: pixelout<=1'b1;
34531: pixelout<=1'b1;
34532: pixelout<=1'b1;
34533: pixelout<=1'b1;
34534: pixelout<=1'b1;
34535: pixelout<=1'b1;
34536: pixelout<=1'b1;
34537: pixelout<=1'b1;
34538: pixelout<=1'b1;
34539: pixelout<=1'b1;
34540: pixelout<=1'b1;
34541: pixelout<=1'b1;
34542: pixelout<=1'b1;
34543: pixelout<=1'b1;
34544: pixelout<=1'b1;
34545: pixelout<=1'b1;
34546: pixelout<=1'b1;
34547: pixelout<=1'b1;
34548: pixelout<=1'b1;
34549: pixelout<=1'b1;
34550: pixelout<=1'b1;
34551: pixelout<=1'b1;
34552: pixelout<=1'b1;
34553: pixelout<=1'b1;
34554: pixelout<=1'b1;
34555: pixelout<=1'b1;
34556: pixelout<=1'b1;
34557: pixelout<=1'b1;
34558: pixelout<=1'b1;
34559: pixelout<=1'b1;
34560: pixelout<=1'b1;
34561: pixelout<=1'b1;
34562: pixelout<=1'b1;
34563: pixelout<=1'b1;
34564: pixelout<=1'b1;
34565: pixelout<=1'b1;
34566: pixelout<=1'b1;
34567: pixelout<=1'b1;
34568: pixelout<=1'b1;
34569: pixelout<=1'b1;
34570: pixelout<=1'b1;
34571: pixelout<=1'b1;
34572: pixelout<=1'b1;
34573: pixelout<=1'b1;
34574: pixelout<=1'b1;
34575: pixelout<=1'b1;
34576: pixelout<=1'b1;
34577: pixelout<=1'b1;
34578: pixelout<=1'b1;
34579: pixelout<=1'b1;
34580: pixelout<=1'b1;
34581: pixelout<=1'b1;
34582: pixelout<=1'b1;
34583: pixelout<=1'b1;
34584: pixelout<=1'b1;
34585: pixelout<=1'b1;
34586: pixelout<=1'b1;
34587: pixelout<=1'b1;
34588: pixelout<=1'b1;
34589: pixelout<=1'b1;
34590: pixelout<=1'b1;
34591: pixelout<=1'b1;
34592: pixelout<=1'b1;
34593: pixelout<=1'b1;
34594: pixelout<=1'b1;
34595: pixelout<=1'b1;
34596: pixelout<=1'b1;
34597: pixelout<=1'b1;
34598: pixelout<=1'b1;
34599: pixelout<=1'b1;
34600: pixelout<=1'b1;
34601: pixelout<=1'b1;
34602: pixelout<=1'b1;
34603: pixelout<=1'b1;
34604: pixelout<=1'b1;
34605: pixelout<=1'b1;
34606: pixelout<=1'b1;
34607: pixelout<=1'b1;
34608: pixelout<=1'b1;
34609: pixelout<=1'b1;
34610: pixelout<=1'b1;
34611: pixelout<=1'b1;
34612: pixelout<=1'b1;
34613: pixelout<=1'b1;
34614: pixelout<=1'b1;
34615: pixelout<=1'b1;
34616: pixelout<=1'b1;
34617: pixelout<=1'b1;
34618: pixelout<=1'b1;
34619: pixelout<=1'b1;
34620: pixelout<=1'b1;
34621: pixelout<=1'b1;
34622: pixelout<=1'b1;
34623: pixelout<=1'b1;
34624: pixelout<=1'b1;
34625: pixelout<=1'b1;
34626: pixelout<=1'b1;
34627: pixelout<=1'b1;
34628: pixelout<=1'b1;
34629: pixelout<=1'b1;
34630: pixelout<=1'b1;
34631: pixelout<=1'b1;
34632: pixelout<=1'b1;
34633: pixelout<=1'b1;
34634: pixelout<=1'b1;
34635: pixelout<=1'b1;
34636: pixelout<=1'b1;
34637: pixelout<=1'b1;
34638: pixelout<=1'b1;
34639: pixelout<=1'b1;
34640: pixelout<=1'b1;
34641: pixelout<=1'b1;
34642: pixelout<=1'b1;
34643: pixelout<=1'b1;
34644: pixelout<=1'b1;
34645: pixelout<=1'b1;
34646: pixelout<=1'b1;
34647: pixelout<=1'b1;
34648: pixelout<=1'b1;
34649: pixelout<=1'b1;
34650: pixelout<=1'b1;
34651: pixelout<=1'b1;
34652: pixelout<=1'b1;
34653: pixelout<=1'b1;
34654: pixelout<=1'b1;
34655: pixelout<=1'b1;
34656: pixelout<=1'b1;
34657: pixelout<=1'b1;
34658: pixelout<=1'b1;
34659: pixelout<=1'b1;
34660: pixelout<=1'b1;
34661: pixelout<=1'b1;
34662: pixelout<=1'b1;
34663: pixelout<=1'b1;
34664: pixelout<=1'b1;
34665: pixelout<=1'b1;
34666: pixelout<=1'b1;
34667: pixelout<=1'b1;
34668: pixelout<=1'b1;
34669: pixelout<=1'b1;
34670: pixelout<=1'b1;
34671: pixelout<=1'b1;
34672: pixelout<=1'b1;
34673: pixelout<=1'b1;
34674: pixelout<=1'b1;
34675: pixelout<=1'b1;
34676: pixelout<=1'b1;
34677: pixelout<=1'b1;
34678: pixelout<=1'b1;
34679: pixelout<=1'b1;
34680: pixelout<=1'b1;
34681: pixelout<=1'b1;
34682: pixelout<=1'b1;
34683: pixelout<=1'b1;
34684: pixelout<=1'b1;
34685: pixelout<=1'b1;
34686: pixelout<=1'b1;
34687: pixelout<=1'b1;
34688: pixelout<=1'b1;
34689: pixelout<=1'b1;
34690: pixelout<=1'b1;
34691: pixelout<=1'b1;
34692: pixelout<=1'b1;
34693: pixelout<=1'b1;
34694: pixelout<=1'b1;
34695: pixelout<=1'b1;
34696: pixelout<=1'b1;
34697: pixelout<=1'b1;
34698: pixelout<=1'b1;
34699: pixelout<=1'b1;
34700: pixelout<=1'b1;
34701: pixelout<=1'b1;
34702: pixelout<=1'b1;
34703: pixelout<=1'b1;
34704: pixelout<=1'b1;
34705: pixelout<=1'b1;
34706: pixelout<=1'b1;
34707: pixelout<=1'b1;
34708: pixelout<=1'b1;
34709: pixelout<=1'b1;
34710: pixelout<=1'b1;
34711: pixelout<=1'b1;
34712: pixelout<=1'b1;
34713: pixelout<=1'b1;
34714: pixelout<=1'b1;
34715: pixelout<=1'b1;
34716: pixelout<=1'b1;
34717: pixelout<=1'b1;
34718: pixelout<=1'b1;
34719: pixelout<=1'b1;
34720: pixelout<=1'b1;
34721: pixelout<=1'b1;
34722: pixelout<=1'b1;
34723: pixelout<=1'b1;
34724: pixelout<=1'b1;
34725: pixelout<=1'b1;
34726: pixelout<=1'b1;
34727: pixelout<=1'b1;
34728: pixelout<=1'b1;
34729: pixelout<=1'b1;
34730: pixelout<=1'b1;
34731: pixelout<=1'b1;
34732: pixelout<=1'b1;
34733: pixelout<=1'b1;
34734: pixelout<=1'b1;
34735: pixelout<=1'b1;
34736: pixelout<=1'b1;
34737: pixelout<=1'b1;
34738: pixelout<=1'b1;
34739: pixelout<=1'b1;
34740: pixelout<=1'b1;
34741: pixelout<=1'b1;
34742: pixelout<=1'b1;
34743: pixelout<=1'b1;
34744: pixelout<=1'b1;
34745: pixelout<=1'b1;
34746: pixelout<=1'b1;
34747: pixelout<=1'b1;
34748: pixelout<=1'b1;
34749: pixelout<=1'b1;
34750: pixelout<=1'b1;
34751: pixelout<=1'b1;
34752: pixelout<=1'b1;
34753: pixelout<=1'b1;
34754: pixelout<=1'b1;
34755: pixelout<=1'b1;
34756: pixelout<=1'b1;
34757: pixelout<=1'b1;
34758: pixelout<=1'b1;
34759: pixelout<=1'b1;
34760: pixelout<=1'b1;
34761: pixelout<=1'b1;
34762: pixelout<=1'b1;
34763: pixelout<=1'b1;
34764: pixelout<=1'b1;
34765: pixelout<=1'b1;
34766: pixelout<=1'b1;
34767: pixelout<=1'b1;
34768: pixelout<=1'b1;
34769: pixelout<=1'b1;
34770: pixelout<=1'b1;
34771: pixelout<=1'b1;
34772: pixelout<=1'b1;
34773: pixelout<=1'b1;
34774: pixelout<=1'b1;
34775: pixelout<=1'b1;
34776: pixelout<=1'b1;
34777: pixelout<=1'b1;
34778: pixelout<=1'b1;
34779: pixelout<=1'b1;
34780: pixelout<=1'b1;
34781: pixelout<=1'b1;
34782: pixelout<=1'b1;
34783: pixelout<=1'b1;
34784: pixelout<=1'b1;
34785: pixelout<=1'b1;
34786: pixelout<=1'b1;
34787: pixelout<=1'b1;
34788: pixelout<=1'b1;
34789: pixelout<=1'b1;
34790: pixelout<=1'b1;
34791: pixelout<=1'b1;
34792: pixelout<=1'b1;
34793: pixelout<=1'b1;
34794: pixelout<=1'b1;
34795: pixelout<=1'b1;
34796: pixelout<=1'b1;
34797: pixelout<=1'b1;
34798: pixelout<=1'b1;
34799: pixelout<=1'b1;
34800: pixelout<=1'b1;
34801: pixelout<=1'b1;
34802: pixelout<=1'b1;
34803: pixelout<=1'b1;
34804: pixelout<=1'b1;
34805: pixelout<=1'b1;
34806: pixelout<=1'b1;
34807: pixelout<=1'b1;
34808: pixelout<=1'b1;
34809: pixelout<=1'b1;
34810: pixelout<=1'b1;
34811: pixelout<=1'b1;
34812: pixelout<=1'b1;
34813: pixelout<=1'b1;
34814: pixelout<=1'b1;
34815: pixelout<=1'b1;
34816: pixelout<=1'b1;
34817: pixelout<=1'b1;
34818: pixelout<=1'b1;
34819: pixelout<=1'b1;
34820: pixelout<=1'b1;
34821: pixelout<=1'b1;
34822: pixelout<=1'b1;
34823: pixelout<=1'b1;
34824: pixelout<=1'b1;
34825: pixelout<=1'b1;
34826: pixelout<=1'b1;
34827: pixelout<=1'b1;
34828: pixelout<=1'b1;
34829: pixelout<=1'b1;
34830: pixelout<=1'b1;
34831: pixelout<=1'b1;
34832: pixelout<=1'b1;
34833: pixelout<=1'b1;
34834: pixelout<=1'b1;
34835: pixelout<=1'b1;
34836: pixelout<=1'b1;
34837: pixelout<=1'b1;
34838: pixelout<=1'b1;
34839: pixelout<=1'b1;
34840: pixelout<=1'b1;
34841: pixelout<=1'b1;
34842: pixelout<=1'b1;
34843: pixelout<=1'b1;
34844: pixelout<=1'b1;
34845: pixelout<=1'b1;
34846: pixelout<=1'b1;
34847: pixelout<=1'b1;
34848: pixelout<=1'b1;
34849: pixelout<=1'b1;
34850: pixelout<=1'b1;
34851: pixelout<=1'b1;
34852: pixelout<=1'b1;
34853: pixelout<=1'b1;
34854: pixelout<=1'b1;
34855: pixelout<=1'b1;
34856: pixelout<=1'b1;
34857: pixelout<=1'b1;
34858: pixelout<=1'b1;
34859: pixelout<=1'b1;
34860: pixelout<=1'b1;
34861: pixelout<=1'b1;
34862: pixelout<=1'b1;
34863: pixelout<=1'b1;
34864: pixelout<=1'b1;
34865: pixelout<=1'b1;
34866: pixelout<=1'b1;
34867: pixelout<=1'b1;
34868: pixelout<=1'b1;
34869: pixelout<=1'b1;
34870: pixelout<=1'b1;
34871: pixelout<=1'b1;
34872: pixelout<=1'b1;
34873: pixelout<=1'b1;
34874: pixelout<=1'b1;
34875: pixelout<=1'b1;
34876: pixelout<=1'b1;
34877: pixelout<=1'b1;
34878: pixelout<=1'b1;
34879: pixelout<=1'b1;
34880: pixelout<=1'b1;
34881: pixelout<=1'b1;
34882: pixelout<=1'b1;
34883: pixelout<=1'b1;
34884: pixelout<=1'b1;
34885: pixelout<=1'b1;
34886: pixelout<=1'b1;
34887: pixelout<=1'b1;
34888: pixelout<=1'b1;
34889: pixelout<=1'b1;
34890: pixelout<=1'b1;
34891: pixelout<=1'b1;
34892: pixelout<=1'b1;
34893: pixelout<=1'b1;
34894: pixelout<=1'b1;
34895: pixelout<=1'b1;
34896: pixelout<=1'b1;
34897: pixelout<=1'b1;
34898: pixelout<=1'b1;
34899: pixelout<=1'b1;
34900: pixelout<=1'b1;
34901: pixelout<=1'b1;
34902: pixelout<=1'b1;
34903: pixelout<=1'b1;
34904: pixelout<=1'b1;
34905: pixelout<=1'b1;
34906: pixelout<=1'b1;
34907: pixelout<=1'b1;
34908: pixelout<=1'b1;
34909: pixelout<=1'b1;
34910: pixelout<=1'b1;
34911: pixelout<=1'b1;
34912: pixelout<=1'b1;
34913: pixelout<=1'b1;
34914: pixelout<=1'b1;
34915: pixelout<=1'b1;
34916: pixelout<=1'b1;
34917: pixelout<=1'b1;
34918: pixelout<=1'b1;
34919: pixelout<=1'b1;
34920: pixelout<=1'b1;
34921: pixelout<=1'b1;
34922: pixelout<=1'b1;
34923: pixelout<=1'b1;
34924: pixelout<=1'b1;
34925: pixelout<=1'b1;
34926: pixelout<=1'b1;
34927: pixelout<=1'b1;
34928: pixelout<=1'b1;
34929: pixelout<=1'b1;
34930: pixelout<=1'b1;
34931: pixelout<=1'b1;
34932: pixelout<=1'b1;
34933: pixelout<=1'b1;
34934: pixelout<=1'b1;
34935: pixelout<=1'b1;
34936: pixelout<=1'b1;
34937: pixelout<=1'b1;
34938: pixelout<=1'b1;
34939: pixelout<=1'b1;
34940: pixelout<=1'b1;
34941: pixelout<=1'b1;
34942: pixelout<=1'b1;
34943: pixelout<=1'b1;
34944: pixelout<=1'b1;
34945: pixelout<=1'b1;
34946: pixelout<=1'b1;
34947: pixelout<=1'b1;
34948: pixelout<=1'b1;
34949: pixelout<=1'b1;
34950: pixelout<=1'b1;
34951: pixelout<=1'b1;
34952: pixelout<=1'b1;
34953: pixelout<=1'b1;
34954: pixelout<=1'b1;
34955: pixelout<=1'b1;
34956: pixelout<=1'b1;
34957: pixelout<=1'b1;
34958: pixelout<=1'b1;
34959: pixelout<=1'b1;
34960: pixelout<=1'b1;
34961: pixelout<=1'b1;
34962: pixelout<=1'b1;
34963: pixelout<=1'b1;
34964: pixelout<=1'b1;
34965: pixelout<=1'b1;
34966: pixelout<=1'b1;
34967: pixelout<=1'b1;
34968: pixelout<=1'b1;
34969: pixelout<=1'b1;
34970: pixelout<=1'b1;
34971: pixelout<=1'b1;
34972: pixelout<=1'b1;
34973: pixelout<=1'b1;
34974: pixelout<=1'b1;
34975: pixelout<=1'b1;
34976: pixelout<=1'b1;
34977: pixelout<=1'b1;
34978: pixelout<=1'b1;
34979: pixelout<=1'b1;
34980: pixelout<=1'b1;
34981: pixelout<=1'b1;
34982: pixelout<=1'b1;
34983: pixelout<=1'b1;
34984: pixelout<=1'b1;
34985: pixelout<=1'b1;
34986: pixelout<=1'b1;
34987: pixelout<=1'b1;
34988: pixelout<=1'b1;
34989: pixelout<=1'b1;
34990: pixelout<=1'b1;
34991: pixelout<=1'b1;
34992: pixelout<=1'b1;
34993: pixelout<=1'b1;
34994: pixelout<=1'b1;
34995: pixelout<=1'b1;
34996: pixelout<=1'b1;
34997: pixelout<=1'b1;
34998: pixelout<=1'b1;
34999: pixelout<=1'b1;
35000: pixelout<=1'b1;
35001: pixelout<=1'b1;
35002: pixelout<=1'b1;
35003: pixelout<=1'b1;
35004: pixelout<=1'b1;
35005: pixelout<=1'b1;
35006: pixelout<=1'b1;
35007: pixelout<=1'b1;
35008: pixelout<=1'b1;
35009: pixelout<=1'b1;
35010: pixelout<=1'b1;
35011: pixelout<=1'b1;
35012: pixelout<=1'b1;
35013: pixelout<=1'b1;
35014: pixelout<=1'b1;
35015: pixelout<=1'b1;
35016: pixelout<=1'b1;
35017: pixelout<=1'b1;
35018: pixelout<=1'b1;
35019: pixelout<=1'b1;
35020: pixelout<=1'b1;
35021: pixelout<=1'b1;
35022: pixelout<=1'b1;
35023: pixelout<=1'b1;
35024: pixelout<=1'b1;
35025: pixelout<=1'b1;
35026: pixelout<=1'b1;
35027: pixelout<=1'b1;
35028: pixelout<=1'b1;
35029: pixelout<=1'b1;
35030: pixelout<=1'b1;
35031: pixelout<=1'b1;
35032: pixelout<=1'b1;
35033: pixelout<=1'b1;
35034: pixelout<=1'b1;
35035: pixelout<=1'b1;
35036: pixelout<=1'b1;
35037: pixelout<=1'b1;
35038: pixelout<=1'b1;
35039: pixelout<=1'b1;
35040: pixelout<=1'b1;
35041: pixelout<=1'b1;
35042: pixelout<=1'b1;
35043: pixelout<=1'b1;
35044: pixelout<=1'b1;
35045: pixelout<=1'b1;
35046: pixelout<=1'b1;
35047: pixelout<=1'b1;
35048: pixelout<=1'b1;
35049: pixelout<=1'b1;
35050: pixelout<=1'b1;
35051: pixelout<=1'b1;
35052: pixelout<=1'b1;
35053: pixelout<=1'b1;
35054: pixelout<=1'b1;
35055: pixelout<=1'b1;
35056: pixelout<=1'b1;
35057: pixelout<=1'b1;
35058: pixelout<=1'b1;
35059: pixelout<=1'b1;
35060: pixelout<=1'b1;
35061: pixelout<=1'b1;
35062: pixelout<=1'b1;
35063: pixelout<=1'b1;
35064: pixelout<=1'b1;
35065: pixelout<=1'b1;
35066: pixelout<=1'b1;
35067: pixelout<=1'b1;
35068: pixelout<=1'b1;
35069: pixelout<=1'b1;
35070: pixelout<=1'b1;
35071: pixelout<=1'b1;
35072: pixelout<=1'b1;
35073: pixelout<=1'b1;
35074: pixelout<=1'b1;
35075: pixelout<=1'b1;
35076: pixelout<=1'b1;
35077: pixelout<=1'b1;
35078: pixelout<=1'b1;
35079: pixelout<=1'b1;
35080: pixelout<=1'b1;
35081: pixelout<=1'b1;
35082: pixelout<=1'b1;
35083: pixelout<=1'b1;
35084: pixelout<=1'b1;
35085: pixelout<=1'b1;
35086: pixelout<=1'b1;
35087: pixelout<=1'b1;
35088: pixelout<=1'b1;
35089: pixelout<=1'b1;
35090: pixelout<=1'b1;
35091: pixelout<=1'b1;
35092: pixelout<=1'b1;
35093: pixelout<=1'b1;
35094: pixelout<=1'b1;
35095: pixelout<=1'b1;
35096: pixelout<=1'b1;
35097: pixelout<=1'b1;
35098: pixelout<=1'b1;
35099: pixelout<=1'b1;
35100: pixelout<=1'b1;
35101: pixelout<=1'b1;
35102: pixelout<=1'b1;
35103: pixelout<=1'b1;
35104: pixelout<=1'b1;
35105: pixelout<=1'b1;
35106: pixelout<=1'b1;
35107: pixelout<=1'b1;
35108: pixelout<=1'b1;
35109: pixelout<=1'b1;
35110: pixelout<=1'b1;
35111: pixelout<=1'b1;
35112: pixelout<=1'b1;
35113: pixelout<=1'b1;
35114: pixelout<=1'b1;
35115: pixelout<=1'b1;
35116: pixelout<=1'b1;
35117: pixelout<=1'b1;
35118: pixelout<=1'b1;
35119: pixelout<=1'b1;
35120: pixelout<=1'b1;
35121: pixelout<=1'b1;
35122: pixelout<=1'b1;
35123: pixelout<=1'b1;
35124: pixelout<=1'b1;
35125: pixelout<=1'b1;
35126: pixelout<=1'b1;
35127: pixelout<=1'b1;
35128: pixelout<=1'b1;
35129: pixelout<=1'b1;
35130: pixelout<=1'b1;
35131: pixelout<=1'b1;
35132: pixelout<=1'b1;
35133: pixelout<=1'b1;
35134: pixelout<=1'b1;
35135: pixelout<=1'b1;
35136: pixelout<=1'b1;
35137: pixelout<=1'b1;
35138: pixelout<=1'b1;
35139: pixelout<=1'b1;
35140: pixelout<=1'b1;
35141: pixelout<=1'b1;
35142: pixelout<=1'b1;
35143: pixelout<=1'b1;
35144: pixelout<=1'b1;
35145: pixelout<=1'b1;
35146: pixelout<=1'b1;
35147: pixelout<=1'b1;
35148: pixelout<=1'b1;
35149: pixelout<=1'b1;
35150: pixelout<=1'b1;
35151: pixelout<=1'b1;
35152: pixelout<=1'b1;
35153: pixelout<=1'b1;
35154: pixelout<=1'b1;
35155: pixelout<=1'b1;
35156: pixelout<=1'b1;
35157: pixelout<=1'b1;
35158: pixelout<=1'b1;
35159: pixelout<=1'b1;
35160: pixelout<=1'b1;
35161: pixelout<=1'b1;
35162: pixelout<=1'b1;
35163: pixelout<=1'b1;
35164: pixelout<=1'b1;
35165: pixelout<=1'b1;
35166: pixelout<=1'b1;
35167: pixelout<=1'b1;
35168: pixelout<=1'b1;
35169: pixelout<=1'b1;
35170: pixelout<=1'b1;
35171: pixelout<=1'b1;
35172: pixelout<=1'b1;
35173: pixelout<=1'b1;
35174: pixelout<=1'b1;
35175: pixelout<=1'b1;
35176: pixelout<=1'b1;
35177: pixelout<=1'b1;
35178: pixelout<=1'b1;
35179: pixelout<=1'b1;
35180: pixelout<=1'b1;
35181: pixelout<=1'b1;
35182: pixelout<=1'b1;
35183: pixelout<=1'b1;
35184: pixelout<=1'b1;
35185: pixelout<=1'b1;
35186: pixelout<=1'b1;
35187: pixelout<=1'b1;
35188: pixelout<=1'b1;
35189: pixelout<=1'b1;
35190: pixelout<=1'b1;
35191: pixelout<=1'b1;
35192: pixelout<=1'b1;
35193: pixelout<=1'b1;
35194: pixelout<=1'b1;
35195: pixelout<=1'b1;
35196: pixelout<=1'b1;
35197: pixelout<=1'b1;
35198: pixelout<=1'b1;
35199: pixelout<=1'b1;
35200: pixelout<=1'b1;
35201: pixelout<=1'b1;
35202: pixelout<=1'b1;
35203: pixelout<=1'b1;
35204: pixelout<=1'b1;
35205: pixelout<=1'b1;
35206: pixelout<=1'b1;
35207: pixelout<=1'b1;
35208: pixelout<=1'b1;
35209: pixelout<=1'b1;
35210: pixelout<=1'b1;
35211: pixelout<=1'b1;
35212: pixelout<=1'b1;
35213: pixelout<=1'b1;
35214: pixelout<=1'b1;
35215: pixelout<=1'b1;
35216: pixelout<=1'b1;
35217: pixelout<=1'b1;
35218: pixelout<=1'b1;
35219: pixelout<=1'b1;
35220: pixelout<=1'b1;
35221: pixelout<=1'b1;
35222: pixelout<=1'b1;
35223: pixelout<=1'b1;
35224: pixelout<=1'b1;
35225: pixelout<=1'b1;
35226: pixelout<=1'b1;
35227: pixelout<=1'b1;
35228: pixelout<=1'b1;
35229: pixelout<=1'b1;
35230: pixelout<=1'b1;
35231: pixelout<=1'b1;
35232: pixelout<=1'b1;
35233: pixelout<=1'b1;
35234: pixelout<=1'b1;
35235: pixelout<=1'b1;
35236: pixelout<=1'b1;
35237: pixelout<=1'b1;
35238: pixelout<=1'b1;
35239: pixelout<=1'b1;
35240: pixelout<=1'b1;
35241: pixelout<=1'b1;
35242: pixelout<=1'b1;
35243: pixelout<=1'b1;
35244: pixelout<=1'b1;
35245: pixelout<=1'b1;
35246: pixelout<=1'b1;
35247: pixelout<=1'b1;
35248: pixelout<=1'b1;
35249: pixelout<=1'b1;
35250: pixelout<=1'b1;
35251: pixelout<=1'b1;
35252: pixelout<=1'b1;
35253: pixelout<=1'b1;
35254: pixelout<=1'b1;
35255: pixelout<=1'b1;
35256: pixelout<=1'b1;
35257: pixelout<=1'b1;
35258: pixelout<=1'b1;
35259: pixelout<=1'b1;
35260: pixelout<=1'b1;
35261: pixelout<=1'b1;
35262: pixelout<=1'b1;
35263: pixelout<=1'b1;
35264: pixelout<=1'b1;
35265: pixelout<=1'b1;
35266: pixelout<=1'b1;
35267: pixelout<=1'b1;
35268: pixelout<=1'b1;
35269: pixelout<=1'b1;
35270: pixelout<=1'b1;
35271: pixelout<=1'b1;
35272: pixelout<=1'b1;
35273: pixelout<=1'b1;
35274: pixelout<=1'b1;
35275: pixelout<=1'b1;
35276: pixelout<=1'b1;
35277: pixelout<=1'b1;
35278: pixelout<=1'b1;
35279: pixelout<=1'b1;
35280: pixelout<=1'b1;
35281: pixelout<=1'b1;
35282: pixelout<=1'b1;
35283: pixelout<=1'b1;
35284: pixelout<=1'b1;
35285: pixelout<=1'b1;
35286: pixelout<=1'b1;
35287: pixelout<=1'b1;
35288: pixelout<=1'b1;
35289: pixelout<=1'b1;
35290: pixelout<=1'b1;
35291: pixelout<=1'b1;
35292: pixelout<=1'b1;
35293: pixelout<=1'b1;
35294: pixelout<=1'b1;
35295: pixelout<=1'b1;
35296: pixelout<=1'b1;
35297: pixelout<=1'b1;
35298: pixelout<=1'b1;
35299: pixelout<=1'b1;
35300: pixelout<=1'b1;
35301: pixelout<=1'b1;
35302: pixelout<=1'b1;
35303: pixelout<=1'b1;
35304: pixelout<=1'b1;
35305: pixelout<=1'b1;
35306: pixelout<=1'b1;
35307: pixelout<=1'b1;
35308: pixelout<=1'b1;
35309: pixelout<=1'b1;
35310: pixelout<=1'b1;
35311: pixelout<=1'b1;
35312: pixelout<=1'b1;
35313: pixelout<=1'b1;
35314: pixelout<=1'b1;
35315: pixelout<=1'b1;
35316: pixelout<=1'b1;
35317: pixelout<=1'b1;
35318: pixelout<=1'b1;
35319: pixelout<=1'b1;
35320: pixelout<=1'b1;
35321: pixelout<=1'b1;
35322: pixelout<=1'b1;
35323: pixelout<=1'b1;
35324: pixelout<=1'b1;
35325: pixelout<=1'b1;
35326: pixelout<=1'b1;
35327: pixelout<=1'b1;
35328: pixelout<=1'b1;
35329: pixelout<=1'b1;
35330: pixelout<=1'b0;
35331: pixelout<=1'b0;
35332: pixelout<=1'b1;
35333: pixelout<=1'b1;
35334: pixelout<=1'b0;
35335: pixelout<=1'b0;
35336: pixelout<=1'b0;
35337: pixelout<=1'b1;
35338: pixelout<=1'b1;
35339: pixelout<=1'b0;
35340: pixelout<=1'b1;
35341: pixelout<=1'b1;
35342: pixelout<=1'b1;
35343: pixelout<=1'b1;
35344: pixelout<=1'b1;
35345: pixelout<=1'b1;
35346: pixelout<=1'b1;
35347: pixelout<=1'b1;
35348: pixelout<=1'b1;
35349: pixelout<=1'b1;
35350: pixelout<=1'b1;
35351: pixelout<=1'b1;
35352: pixelout<=1'b1;
35353: pixelout<=1'b1;
35354: pixelout<=1'b1;
35355: pixelout<=1'b1;
35356: pixelout<=1'b1;
35357: pixelout<=1'b1;
35358: pixelout<=1'b1;
35359: pixelout<=1'b1;
35360: pixelout<=1'b1;
35361: pixelout<=1'b1;
35362: pixelout<=1'b1;
35363: pixelout<=1'b1;
35364: pixelout<=1'b1;
35365: pixelout<=1'b1;
35366: pixelout<=1'b1;
35367: pixelout<=1'b1;
35368: pixelout<=1'b1;
35369: pixelout<=1'b1;
35370: pixelout<=1'b1;
35371: pixelout<=1'b1;
35372: pixelout<=1'b1;
35373: pixelout<=1'b1;
35374: pixelout<=1'b1;
35375: pixelout<=1'b1;
35376: pixelout<=1'b1;
35377: pixelout<=1'b1;
35378: pixelout<=1'b1;
35379: pixelout<=1'b1;
35380: pixelout<=1'b1;
35381: pixelout<=1'b1;
35382: pixelout<=1'b1;
35383: pixelout<=1'b1;
35384: pixelout<=1'b1;
35385: pixelout<=1'b1;
35386: pixelout<=1'b1;
35387: pixelout<=1'b1;
35388: pixelout<=1'b1;
35389: pixelout<=1'b1;
35390: pixelout<=1'b1;
35391: pixelout<=1'b1;
35392: pixelout<=1'b1;
35393: pixelout<=1'b1;
35394: pixelout<=1'b1;
35395: pixelout<=1'b1;
35396: pixelout<=1'b1;
35397: pixelout<=1'b1;
35398: pixelout<=1'b1;
35399: pixelout<=1'b1;
35400: pixelout<=1'b1;
35401: pixelout<=1'b1;
35402: pixelout<=1'b1;
35403: pixelout<=1'b1;
35404: pixelout<=1'b1;
35405: pixelout<=1'b1;
35406: pixelout<=1'b1;
35407: pixelout<=1'b1;
35408: pixelout<=1'b1;
35409: pixelout<=1'b1;
35410: pixelout<=1'b1;
35411: pixelout<=1'b1;
35412: pixelout<=1'b1;
35413: pixelout<=1'b1;
35414: pixelout<=1'b1;
35415: pixelout<=1'b1;
35416: pixelout<=1'b1;
35417: pixelout<=1'b1;
35418: pixelout<=1'b1;
35419: pixelout<=1'b1;
35420: pixelout<=1'b1;
35421: pixelout<=1'b1;
35422: pixelout<=1'b1;
35423: pixelout<=1'b1;
35424: pixelout<=1'b1;
35425: pixelout<=1'b1;
35426: pixelout<=1'b1;
35427: pixelout<=1'b1;
35428: pixelout<=1'b1;
35429: pixelout<=1'b1;
35430: pixelout<=1'b1;
35431: pixelout<=1'b1;
35432: pixelout<=1'b1;
35433: pixelout<=1'b1;
35434: pixelout<=1'b1;
35435: pixelout<=1'b1;
35436: pixelout<=1'b1;
35437: pixelout<=1'b1;
35438: pixelout<=1'b1;
35439: pixelout<=1'b1;
35440: pixelout<=1'b1;
35441: pixelout<=1'b1;
35442: pixelout<=1'b1;
35443: pixelout<=1'b1;
35444: pixelout<=1'b1;
35445: pixelout<=1'b1;
35446: pixelout<=1'b1;
35447: pixelout<=1'b1;
35448: pixelout<=1'b1;
35449: pixelout<=1'b1;
35450: pixelout<=1'b1;
35451: pixelout<=1'b1;
35452: pixelout<=1'b1;
35453: pixelout<=1'b1;
35454: pixelout<=1'b1;
35455: pixelout<=1'b1;
35456: pixelout<=1'b1;
35457: pixelout<=1'b1;
35458: pixelout<=1'b1;
35459: pixelout<=1'b1;
35460: pixelout<=1'b1;
35461: pixelout<=1'b1;
35462: pixelout<=1'b1;
35463: pixelout<=1'b1;
35464: pixelout<=1'b1;
35465: pixelout<=1'b1;
35466: pixelout<=1'b1;
35467: pixelout<=1'b1;
35468: pixelout<=1'b1;
35469: pixelout<=1'b1;
35470: pixelout<=1'b1;
35471: pixelout<=1'b1;
35472: pixelout<=1'b1;
35473: pixelout<=1'b1;
35474: pixelout<=1'b1;
35475: pixelout<=1'b1;
35476: pixelout<=1'b1;
35477: pixelout<=1'b1;
35478: pixelout<=1'b1;
35479: pixelout<=1'b1;
35480: pixelout<=1'b1;
35481: pixelout<=1'b1;
35482: pixelout<=1'b1;
35483: pixelout<=1'b1;
35484: pixelout<=1'b1;
35485: pixelout<=1'b1;
35486: pixelout<=1'b1;
35487: pixelout<=1'b1;
35488: pixelout<=1'b1;
35489: pixelout<=1'b1;
35490: pixelout<=1'b1;
35491: pixelout<=1'b1;
35492: pixelout<=1'b1;
35493: pixelout<=1'b1;
35494: pixelout<=1'b1;
35495: pixelout<=1'b1;
35496: pixelout<=1'b1;
35497: pixelout<=1'b1;
35498: pixelout<=1'b1;
35499: pixelout<=1'b1;
35500: pixelout<=1'b1;
35501: pixelout<=1'b1;
35502: pixelout<=1'b1;
35503: pixelout<=1'b1;
35504: pixelout<=1'b1;
35505: pixelout<=1'b1;
35506: pixelout<=1'b1;
35507: pixelout<=1'b1;
35508: pixelout<=1'b1;
35509: pixelout<=1'b1;
35510: pixelout<=1'b1;
35511: pixelout<=1'b1;
35512: pixelout<=1'b1;
35513: pixelout<=1'b1;
35514: pixelout<=1'b1;
35515: pixelout<=1'b1;
35516: pixelout<=1'b1;
35517: pixelout<=1'b1;
35518: pixelout<=1'b1;
35519: pixelout<=1'b1;
35520: pixelout<=1'b1;
35521: pixelout<=1'b1;
35522: pixelout<=1'b1;
35523: pixelout<=1'b1;
35524: pixelout<=1'b1;
35525: pixelout<=1'b1;
35526: pixelout<=1'b1;
35527: pixelout<=1'b1;
35528: pixelout<=1'b1;
35529: pixelout<=1'b1;
35530: pixelout<=1'b1;
35531: pixelout<=1'b1;
35532: pixelout<=1'b1;
35533: pixelout<=1'b1;
35534: pixelout<=1'b1;
35535: pixelout<=1'b1;
35536: pixelout<=1'b1;
35537: pixelout<=1'b1;
35538: pixelout<=1'b1;
35539: pixelout<=1'b1;
35540: pixelout<=1'b1;
35541: pixelout<=1'b1;
35542: pixelout<=1'b1;
35543: pixelout<=1'b1;
35544: pixelout<=1'b1;
35545: pixelout<=1'b0;
35546: pixelout<=1'b1;
35547: pixelout<=1'b1;
35548: pixelout<=1'b1;
35549: pixelout<=1'b1;
35550: pixelout<=1'b1;
35551: pixelout<=1'b1;
35552: pixelout<=1'b1;
35553: pixelout<=1'b1;
35554: pixelout<=1'b1;
35555: pixelout<=1'b1;
35556: pixelout<=1'b0;
35557: pixelout<=1'b1;
35558: pixelout<=1'b1;
35559: pixelout<=1'b1;
35560: pixelout<=1'b1;
35561: pixelout<=1'b1;
35562: pixelout<=1'b1;
35563: pixelout<=1'b1;
35564: pixelout<=1'b1;
35565: pixelout<=1'b1;
35566: pixelout<=1'b1;
35567: pixelout<=1'b1;
35568: pixelout<=1'b1;
35569: pixelout<=1'b1;
35570: pixelout<=1'b1;
35571: pixelout<=1'b1;
35572: pixelout<=1'b0;
35573: pixelout<=1'b1;
35574: pixelout<=1'b1;
35575: pixelout<=1'b1;
35576: pixelout<=1'b1;
35577: pixelout<=1'b1;
35578: pixelout<=1'b1;
35579: pixelout<=1'b0;
35580: pixelout<=1'b1;
35581: pixelout<=1'b1;
35582: pixelout<=1'b1;
35583: pixelout<=1'b1;
35584: pixelout<=1'b1;
35585: pixelout<=1'b1;
35586: pixelout<=1'b1;
35587: pixelout<=1'b1;
35588: pixelout<=1'b1;
35589: pixelout<=1'b1;
35590: pixelout<=1'b1;
35591: pixelout<=1'b1;
35592: pixelout<=1'b1;
35593: pixelout<=1'b1;
35594: pixelout<=1'b1;
35595: pixelout<=1'b1;
35596: pixelout<=1'b1;
35597: pixelout<=1'b1;
35598: pixelout<=1'b1;
35599: pixelout<=1'b1;
35600: pixelout<=1'b1;
35601: pixelout<=1'b1;
35602: pixelout<=1'b1;
35603: pixelout<=1'b1;
35604: pixelout<=1'b1;
35605: pixelout<=1'b1;
35606: pixelout<=1'b1;
35607: pixelout<=1'b1;
35608: pixelout<=1'b1;
35609: pixelout<=1'b1;
35610: pixelout<=1'b1;
35611: pixelout<=1'b1;
35612: pixelout<=1'b1;
35613: pixelout<=1'b1;
35614: pixelout<=1'b1;
35615: pixelout<=1'b1;
35616: pixelout<=1'b1;
35617: pixelout<=1'b1;
35618: pixelout<=1'b1;
35619: pixelout<=1'b1;
35620: pixelout<=1'b1;
35621: pixelout<=1'b1;
35622: pixelout<=1'b1;
35623: pixelout<=1'b1;
35624: pixelout<=1'b1;
35625: pixelout<=1'b1;
35626: pixelout<=1'b1;
35627: pixelout<=1'b1;
35628: pixelout<=1'b1;
35629: pixelout<=1'b1;
35630: pixelout<=1'b1;
35631: pixelout<=1'b1;
35632: pixelout<=1'b1;
35633: pixelout<=1'b1;
35634: pixelout<=1'b1;
35635: pixelout<=1'b1;
35636: pixelout<=1'b1;
35637: pixelout<=1'b1;
35638: pixelout<=1'b1;
35639: pixelout<=1'b1;
35640: pixelout<=1'b1;
35641: pixelout<=1'b1;
35642: pixelout<=1'b1;
35643: pixelout<=1'b1;
35644: pixelout<=1'b1;
35645: pixelout<=1'b1;
35646: pixelout<=1'b1;
35647: pixelout<=1'b1;
35648: pixelout<=1'b1;
35649: pixelout<=1'b1;
35650: pixelout<=1'b1;
35651: pixelout<=1'b1;
35652: pixelout<=1'b1;
35653: pixelout<=1'b1;
35654: pixelout<=1'b1;
35655: pixelout<=1'b1;
35656: pixelout<=1'b1;
35657: pixelout<=1'b1;
35658: pixelout<=1'b1;
35659: pixelout<=1'b1;
35660: pixelout<=1'b1;
35661: pixelout<=1'b1;
35662: pixelout<=1'b1;
35663: pixelout<=1'b1;
35664: pixelout<=1'b1;
35665: pixelout<=1'b1;
35666: pixelout<=1'b1;
35667: pixelout<=1'b1;
35668: pixelout<=1'b1;
35669: pixelout<=1'b1;
35670: pixelout<=1'b1;
35671: pixelout<=1'b1;
35672: pixelout<=1'b1;
35673: pixelout<=1'b1;
35674: pixelout<=1'b1;
35675: pixelout<=1'b1;
35676: pixelout<=1'b1;
35677: pixelout<=1'b1;
35678: pixelout<=1'b1;
35679: pixelout<=1'b1;
35680: pixelout<=1'b1;
35681: pixelout<=1'b1;
35682: pixelout<=1'b1;
35683: pixelout<=1'b1;
35684: pixelout<=1'b1;
35685: pixelout<=1'b1;
35686: pixelout<=1'b1;
35687: pixelout<=1'b1;
35688: pixelout<=1'b1;
35689: pixelout<=1'b1;
35690: pixelout<=1'b1;
35691: pixelout<=1'b1;
35692: pixelout<=1'b1;
35693: pixelout<=1'b1;
35694: pixelout<=1'b1;
35695: pixelout<=1'b1;
35696: pixelout<=1'b1;
35697: pixelout<=1'b1;
35698: pixelout<=1'b1;
35699: pixelout<=1'b1;
35700: pixelout<=1'b1;
35701: pixelout<=1'b1;
35702: pixelout<=1'b1;
35703: pixelout<=1'b1;
35704: pixelout<=1'b1;
35705: pixelout<=1'b1;
35706: pixelout<=1'b1;
35707: pixelout<=1'b1;
35708: pixelout<=1'b1;
35709: pixelout<=1'b1;
35710: pixelout<=1'b1;
35711: pixelout<=1'b1;
35712: pixelout<=1'b1;
35713: pixelout<=1'b1;
35714: pixelout<=1'b1;
35715: pixelout<=1'b1;
35716: pixelout<=1'b1;
35717: pixelout<=1'b1;
35718: pixelout<=1'b1;
35719: pixelout<=1'b1;
35720: pixelout<=1'b1;
35721: pixelout<=1'b1;
35722: pixelout<=1'b1;
35723: pixelout<=1'b1;
35724: pixelout<=1'b1;
35725: pixelout<=1'b1;
35726: pixelout<=1'b1;
35727: pixelout<=1'b1;
35728: pixelout<=1'b1;
35729: pixelout<=1'b1;
35730: pixelout<=1'b1;
35731: pixelout<=1'b1;
35732: pixelout<=1'b1;
35733: pixelout<=1'b1;
35734: pixelout<=1'b1;
35735: pixelout<=1'b1;
35736: pixelout<=1'b1;
35737: pixelout<=1'b1;
35738: pixelout<=1'b1;
35739: pixelout<=1'b1;
35740: pixelout<=1'b1;
35741: pixelout<=1'b1;
35742: pixelout<=1'b1;
35743: pixelout<=1'b1;
35744: pixelout<=1'b1;
35745: pixelout<=1'b1;
35746: pixelout<=1'b1;
35747: pixelout<=1'b1;
35748: pixelout<=1'b1;
35749: pixelout<=1'b1;
35750: pixelout<=1'b1;
35751: pixelout<=1'b1;
35752: pixelout<=1'b1;
35753: pixelout<=1'b1;
35754: pixelout<=1'b1;
35755: pixelout<=1'b1;
35756: pixelout<=1'b1;
35757: pixelout<=1'b1;
35758: pixelout<=1'b1;
35759: pixelout<=1'b1;
35760: pixelout<=1'b1;
35761: pixelout<=1'b1;
35762: pixelout<=1'b1;
35763: pixelout<=1'b1;
35764: pixelout<=1'b1;
35765: pixelout<=1'b1;
35766: pixelout<=1'b1;
35767: pixelout<=1'b1;
35768: pixelout<=1'b1;
35769: pixelout<=1'b1;
35770: pixelout<=1'b1;
35771: pixelout<=1'b1;
35772: pixelout<=1'b1;
35773: pixelout<=1'b1;
35774: pixelout<=1'b1;
35775: pixelout<=1'b1;
35776: pixelout<=1'b1;
35777: pixelout<=1'b1;
35778: pixelout<=1'b1;
35779: pixelout<=1'b1;
35780: pixelout<=1'b1;
35781: pixelout<=1'b1;
35782: pixelout<=1'b1;
35783: pixelout<=1'b1;
35784: pixelout<=1'b1;
35785: pixelout<=1'b1;
35786: pixelout<=1'b1;
35787: pixelout<=1'b1;
35788: pixelout<=1'b1;
35789: pixelout<=1'b1;
35790: pixelout<=1'b1;
35791: pixelout<=1'b1;
35792: pixelout<=1'b1;
35793: pixelout<=1'b1;
35794: pixelout<=1'b1;
35795: pixelout<=1'b1;
35796: pixelout<=1'b0;
35797: pixelout<=1'b1;
35798: pixelout<=1'b1;
35799: pixelout<=1'b1;
35800: pixelout<=1'b1;
35801: pixelout<=1'b1;
35802: pixelout<=1'b1;
35803: pixelout<=1'b1;
35804: pixelout<=1'b1;
35805: pixelout<=1'b1;
35806: pixelout<=1'b1;
35807: pixelout<=1'b1;
35808: pixelout<=1'b1;
35809: pixelout<=1'b1;
35810: pixelout<=1'b1;
35811: pixelout<=1'b1;
35812: pixelout<=1'b0;
35813: pixelout<=1'b1;
35814: pixelout<=1'b1;
35815: pixelout<=1'b1;
35816: pixelout<=1'b1;
35817: pixelout<=1'b1;
35818: pixelout<=1'b1;
35819: pixelout<=1'b0;
35820: pixelout<=1'b1;
35821: pixelout<=1'b1;
35822: pixelout<=1'b1;
35823: pixelout<=1'b0;
35824: pixelout<=1'b1;
35825: pixelout<=1'b1;
35826: pixelout<=1'b1;
35827: pixelout<=1'b1;
35828: pixelout<=1'b1;
35829: pixelout<=1'b1;
35830: pixelout<=1'b0;
35831: pixelout<=1'b1;
35832: pixelout<=1'b1;
35833: pixelout<=1'b1;
35834: pixelout<=1'b1;
35835: pixelout<=1'b1;
35836: pixelout<=1'b1;
35837: pixelout<=1'b1;
35838: pixelout<=1'b1;
35839: pixelout<=1'b1;
35840: pixelout<=1'b1;
35841: pixelout<=1'b1;
35842: pixelout<=1'b1;
35843: pixelout<=1'b1;
35844: pixelout<=1'b1;
35845: pixelout<=1'b1;
35846: pixelout<=1'b1;
35847: pixelout<=1'b1;
35848: pixelout<=1'b1;
35849: pixelout<=1'b1;
35850: pixelout<=1'b1;
35851: pixelout<=1'b1;
35852: pixelout<=1'b1;
35853: pixelout<=1'b1;
35854: pixelout<=1'b1;
35855: pixelout<=1'b1;
35856: pixelout<=1'b1;
35857: pixelout<=1'b1;
35858: pixelout<=1'b1;
35859: pixelout<=1'b1;
35860: pixelout<=1'b1;
35861: pixelout<=1'b1;
35862: pixelout<=1'b1;
35863: pixelout<=1'b1;
35864: pixelout<=1'b1;
35865: pixelout<=1'b1;
35866: pixelout<=1'b1;
35867: pixelout<=1'b1;
35868: pixelout<=1'b1;
35869: pixelout<=1'b1;
35870: pixelout<=1'b1;
35871: pixelout<=1'b1;
35872: pixelout<=1'b1;
35873: pixelout<=1'b1;
35874: pixelout<=1'b1;
35875: pixelout<=1'b1;
35876: pixelout<=1'b1;
35877: pixelout<=1'b1;
35878: pixelout<=1'b1;
35879: pixelout<=1'b1;
35880: pixelout<=1'b1;
35881: pixelout<=1'b1;
35882: pixelout<=1'b1;
35883: pixelout<=1'b1;
35884: pixelout<=1'b1;
35885: pixelout<=1'b1;
35886: pixelout<=1'b1;
35887: pixelout<=1'b1;
35888: pixelout<=1'b1;
35889: pixelout<=1'b1;
35890: pixelout<=1'b1;
35891: pixelout<=1'b1;
35892: pixelout<=1'b1;
35893: pixelout<=1'b1;
35894: pixelout<=1'b1;
35895: pixelout<=1'b1;
35896: pixelout<=1'b1;
35897: pixelout<=1'b1;
35898: pixelout<=1'b1;
35899: pixelout<=1'b1;
35900: pixelout<=1'b1;
35901: pixelout<=1'b1;
35902: pixelout<=1'b1;
35903: pixelout<=1'b1;
35904: pixelout<=1'b1;
35905: pixelout<=1'b1;
35906: pixelout<=1'b1;
35907: pixelout<=1'b1;
35908: pixelout<=1'b1;
35909: pixelout<=1'b1;
35910: pixelout<=1'b1;
35911: pixelout<=1'b1;
35912: pixelout<=1'b1;
35913: pixelout<=1'b1;
35914: pixelout<=1'b1;
35915: pixelout<=1'b1;
35916: pixelout<=1'b1;
35917: pixelout<=1'b1;
35918: pixelout<=1'b1;
35919: pixelout<=1'b1;
35920: pixelout<=1'b1;
35921: pixelout<=1'b1;
35922: pixelout<=1'b1;
35923: pixelout<=1'b1;
35924: pixelout<=1'b1;
35925: pixelout<=1'b1;
35926: pixelout<=1'b0;
35927: pixelout<=1'b1;
35928: pixelout<=1'b1;
35929: pixelout<=1'b1;
35930: pixelout<=1'b1;
35931: pixelout<=1'b1;
35932: pixelout<=1'b1;
35933: pixelout<=1'b1;
35934: pixelout<=1'b1;
35935: pixelout<=1'b1;
35936: pixelout<=1'b1;
35937: pixelout<=1'b1;
35938: pixelout<=1'b1;
35939: pixelout<=1'b1;
35940: pixelout<=1'b1;
35941: pixelout<=1'b1;
35942: pixelout<=1'b1;
35943: pixelout<=1'b1;
35944: pixelout<=1'b1;
35945: pixelout<=1'b1;
35946: pixelout<=1'b1;
35947: pixelout<=1'b1;
35948: pixelout<=1'b1;
35949: pixelout<=1'b1;
35950: pixelout<=1'b1;
35951: pixelout<=1'b1;
35952: pixelout<=1'b1;
35953: pixelout<=1'b1;
35954: pixelout<=1'b1;
35955: pixelout<=1'b1;
35956: pixelout<=1'b1;
35957: pixelout<=1'b1;
35958: pixelout<=1'b1;
35959: pixelout<=1'b1;
35960: pixelout<=1'b1;
35961: pixelout<=1'b1;
35962: pixelout<=1'b1;
35963: pixelout<=1'b1;
35964: pixelout<=1'b0;
35965: pixelout<=1'b1;
35966: pixelout<=1'b1;
35967: pixelout<=1'b1;
35968: pixelout<=1'b1;
35969: pixelout<=1'b1;
35970: pixelout<=1'b1;
35971: pixelout<=1'b1;
35972: pixelout<=1'b1;
35973: pixelout<=1'b1;
35974: pixelout<=1'b1;
35975: pixelout<=1'b1;
35976: pixelout<=1'b1;
35977: pixelout<=1'b1;
35978: pixelout<=1'b1;
35979: pixelout<=1'b1;
35980: pixelout<=1'b1;
35981: pixelout<=1'b1;
35982: pixelout<=1'b1;
35983: pixelout<=1'b1;
35984: pixelout<=1'b1;
35985: pixelout<=1'b1;
35986: pixelout<=1'b1;
35987: pixelout<=1'b1;
35988: pixelout<=1'b1;
35989: pixelout<=1'b1;
35990: pixelout<=1'b1;
35991: pixelout<=1'b1;
35992: pixelout<=1'b1;
35993: pixelout<=1'b1;
35994: pixelout<=1'b1;
35995: pixelout<=1'b1;
35996: pixelout<=1'b1;
35997: pixelout<=1'b1;
35998: pixelout<=1'b1;
35999: pixelout<=1'b1;
36000: pixelout<=1'b1;
36001: pixelout<=1'b1;
36002: pixelout<=1'b1;
36003: pixelout<=1'b1;
36004: pixelout<=1'b1;
36005: pixelout<=1'b0;
36006: pixelout<=1'b0;
36007: pixelout<=1'b1;
36008: pixelout<=1'b1;
36009: pixelout<=1'b1;
36010: pixelout<=1'b0;
36011: pixelout<=1'b0;
36012: pixelout<=1'b1;
36013: pixelout<=1'b1;
36014: pixelout<=1'b1;
36015: pixelout<=1'b0;
36016: pixelout<=1'b0;
36017: pixelout<=1'b1;
36018: pixelout<=1'b1;
36019: pixelout<=1'b0;
36020: pixelout<=1'b0;
36021: pixelout<=1'b0;
36022: pixelout<=1'b1;
36023: pixelout<=1'b1;
36024: pixelout<=1'b1;
36025: pixelout<=1'b1;
36026: pixelout<=1'b1;
36027: pixelout<=1'b0;
36028: pixelout<=1'b1;
36029: pixelout<=1'b0;
36030: pixelout<=1'b1;
36031: pixelout<=1'b1;
36032: pixelout<=1'b1;
36033: pixelout<=1'b0;
36034: pixelout<=1'b0;
36035: pixelout<=1'b1;
36036: pixelout<=1'b0;
36037: pixelout<=1'b1;
36038: pixelout<=1'b1;
36039: pixelout<=1'b1;
36040: pixelout<=1'b1;
36041: pixelout<=1'b1;
36042: pixelout<=1'b1;
36043: pixelout<=1'b1;
36044: pixelout<=1'b0;
36045: pixelout<=1'b0;
36046: pixelout<=1'b1;
36047: pixelout<=1'b1;
36048: pixelout<=1'b1;
36049: pixelout<=1'b1;
36050: pixelout<=1'b0;
36051: pixelout<=1'b0;
36052: pixelout<=1'b1;
36053: pixelout<=1'b1;
36054: pixelout<=1'b0;
36055: pixelout<=1'b0;
36056: pixelout<=1'b0;
36057: pixelout<=1'b1;
36058: pixelout<=1'b1;
36059: pixelout<=1'b0;
36060: pixelout<=1'b1;
36061: pixelout<=1'b1;
36062: pixelout<=1'b1;
36063: pixelout<=1'b1;
36064: pixelout<=1'b1;
36065: pixelout<=1'b0;
36066: pixelout<=1'b0;
36067: pixelout<=1'b0;
36068: pixelout<=1'b0;
36069: pixelout<=1'b1;
36070: pixelout<=1'b1;
36071: pixelout<=1'b1;
36072: pixelout<=1'b1;
36073: pixelout<=1'b1;
36074: pixelout<=1'b1;
36075: pixelout<=1'b1;
36076: pixelout<=1'b1;
36077: pixelout<=1'b1;
36078: pixelout<=1'b1;
36079: pixelout<=1'b1;
36080: pixelout<=1'b1;
36081: pixelout<=1'b1;
36082: pixelout<=1'b1;
36083: pixelout<=1'b1;
36084: pixelout<=1'b1;
36085: pixelout<=1'b1;
36086: pixelout<=1'b1;
36087: pixelout<=1'b1;
36088: pixelout<=1'b1;
36089: pixelout<=1'b1;
36090: pixelout<=1'b1;
36091: pixelout<=1'b1;
36092: pixelout<=1'b1;
36093: pixelout<=1'b1;
36094: pixelout<=1'b1;
36095: pixelout<=1'b1;
36096: pixelout<=1'b1;
36097: pixelout<=1'b1;
36098: pixelout<=1'b1;
36099: pixelout<=1'b1;
36100: pixelout<=1'b1;
36101: pixelout<=1'b1;
36102: pixelout<=1'b1;
36103: pixelout<=1'b1;
36104: pixelout<=1'b1;
36105: pixelout<=1'b1;
36106: pixelout<=1'b1;
36107: pixelout<=1'b1;
36108: pixelout<=1'b1;
36109: pixelout<=1'b1;
36110: pixelout<=1'b1;
36111: pixelout<=1'b1;
36112: pixelout<=1'b1;
36113: pixelout<=1'b1;
36114: pixelout<=1'b1;
36115: pixelout<=1'b1;
36116: pixelout<=1'b1;
36117: pixelout<=1'b1;
36118: pixelout<=1'b1;
36119: pixelout<=1'b1;
36120: pixelout<=1'b1;
36121: pixelout<=1'b1;
36122: pixelout<=1'b1;
36123: pixelout<=1'b1;
36124: pixelout<=1'b1;
36125: pixelout<=1'b1;
36126: pixelout<=1'b1;
36127: pixelout<=1'b1;
36128: pixelout<=1'b1;
36129: pixelout<=1'b1;
36130: pixelout<=1'b1;
36131: pixelout<=1'b1;
36132: pixelout<=1'b1;
36133: pixelout<=1'b1;
36134: pixelout<=1'b1;
36135: pixelout<=1'b1;
36136: pixelout<=1'b1;
36137: pixelout<=1'b1;
36138: pixelout<=1'b1;
36139: pixelout<=1'b1;
36140: pixelout<=1'b1;
36141: pixelout<=1'b1;
36142: pixelout<=1'b1;
36143: pixelout<=1'b1;
36144: pixelout<=1'b1;
36145: pixelout<=1'b1;
36146: pixelout<=1'b1;
36147: pixelout<=1'b1;
36148: pixelout<=1'b1;
36149: pixelout<=1'b1;
36150: pixelout<=1'b1;
36151: pixelout<=1'b1;
36152: pixelout<=1'b1;
36153: pixelout<=1'b1;
36154: pixelout<=1'b1;
36155: pixelout<=1'b1;
36156: pixelout<=1'b1;
36157: pixelout<=1'b1;
36158: pixelout<=1'b1;
36159: pixelout<=1'b1;
36160: pixelout<=1'b1;
36161: pixelout<=1'b1;
36162: pixelout<=1'b1;
36163: pixelout<=1'b1;
36164: pixelout<=1'b1;
36165: pixelout<=1'b1;
36166: pixelout<=1'b1;
36167: pixelout<=1'b1;
36168: pixelout<=1'b1;
36169: pixelout<=1'b1;
36170: pixelout<=1'b1;
36171: pixelout<=1'b1;
36172: pixelout<=1'b1;
36173: pixelout<=1'b1;
36174: pixelout<=1'b1;
36175: pixelout<=1'b0;
36176: pixelout<=1'b1;
36177: pixelout<=1'b1;
36178: pixelout<=1'b1;
36179: pixelout<=1'b1;
36180: pixelout<=1'b1;
36181: pixelout<=1'b1;
36182: pixelout<=1'b1;
36183: pixelout<=1'b1;
36184: pixelout<=1'b1;
36185: pixelout<=1'b1;
36186: pixelout<=1'b1;
36187: pixelout<=1'b1;
36188: pixelout<=1'b1;
36189: pixelout<=1'b0;
36190: pixelout<=1'b1;
36191: pixelout<=1'b1;
36192: pixelout<=1'b1;
36193: pixelout<=1'b1;
36194: pixelout<=1'b1;
36195: pixelout<=1'b1;
36196: pixelout<=1'b1;
36197: pixelout<=1'b1;
36198: pixelout<=1'b1;
36199: pixelout<=1'b1;
36200: pixelout<=1'b1;
36201: pixelout<=1'b1;
36202: pixelout<=1'b1;
36203: pixelout<=1'b1;
36204: pixelout<=1'b0;
36205: pixelout<=1'b1;
36206: pixelout<=1'b1;
36207: pixelout<=1'b1;
36208: pixelout<=1'b1;
36209: pixelout<=1'b1;
36210: pixelout<=1'b1;
36211: pixelout<=1'b1;
36212: pixelout<=1'b1;
36213: pixelout<=1'b1;
36214: pixelout<=1'b1;
36215: pixelout<=1'b1;
36216: pixelout<=1'b1;
36217: pixelout<=1'b1;
36218: pixelout<=1'b1;
36219: pixelout<=1'b1;
36220: pixelout<=1'b1;
36221: pixelout<=1'b1;
36222: pixelout<=1'b1;
36223: pixelout<=1'b1;
36224: pixelout<=1'b1;
36225: pixelout<=1'b1;
36226: pixelout<=1'b1;
36227: pixelout<=1'b1;
36228: pixelout<=1'b1;
36229: pixelout<=1'b1;
36230: pixelout<=1'b1;
36231: pixelout<=1'b1;
36232: pixelout<=1'b1;
36233: pixelout<=1'b1;
36234: pixelout<=1'b1;
36235: pixelout<=1'b1;
36236: pixelout<=1'b1;
36237: pixelout<=1'b1;
36238: pixelout<=1'b1;
36239: pixelout<=1'b1;
36240: pixelout<=1'b1;
36241: pixelout<=1'b1;
36242: pixelout<=1'b1;
36243: pixelout<=1'b1;
36244: pixelout<=1'b0;
36245: pixelout<=1'b1;
36246: pixelout<=1'b1;
36247: pixelout<=1'b0;
36248: pixelout<=1'b1;
36249: pixelout<=1'b0;
36250: pixelout<=1'b1;
36251: pixelout<=1'b1;
36252: pixelout<=1'b0;
36253: pixelout<=1'b1;
36254: pixelout<=1'b1;
36255: pixelout<=1'b1;
36256: pixelout<=1'b1;
36257: pixelout<=1'b0;
36258: pixelout<=1'b1;
36259: pixelout<=1'b1;
36260: pixelout<=1'b1;
36261: pixelout<=1'b1;
36262: pixelout<=1'b1;
36263: pixelout<=1'b1;
36264: pixelout<=1'b1;
36265: pixelout<=1'b1;
36266: pixelout<=1'b1;
36267: pixelout<=1'b0;
36268: pixelout<=1'b1;
36269: pixelout<=1'b0;
36270: pixelout<=1'b1;
36271: pixelout<=1'b1;
36272: pixelout<=1'b1;
36273: pixelout<=1'b1;
36274: pixelout<=1'b1;
36275: pixelout<=1'b1;
36276: pixelout<=1'b0;
36277: pixelout<=1'b1;
36278: pixelout<=1'b1;
36279: pixelout<=1'b1;
36280: pixelout<=1'b1;
36281: pixelout<=1'b1;
36282: pixelout<=1'b1;
36283: pixelout<=1'b1;
36284: pixelout<=1'b1;
36285: pixelout<=1'b1;
36286: pixelout<=1'b0;
36287: pixelout<=1'b1;
36288: pixelout<=1'b1;
36289: pixelout<=1'b1;
36290: pixelout<=1'b1;
36291: pixelout<=1'b1;
36292: pixelout<=1'b0;
36293: pixelout<=1'b1;
36294: pixelout<=1'b1;
36295: pixelout<=1'b1;
36296: pixelout<=1'b1;
36297: pixelout<=1'b1;
36298: pixelout<=1'b1;
36299: pixelout<=1'b0;
36300: pixelout<=1'b1;
36301: pixelout<=1'b1;
36302: pixelout<=1'b1;
36303: pixelout<=1'b1;
36304: pixelout<=1'b1;
36305: pixelout<=1'b1;
36306: pixelout<=1'b1;
36307: pixelout<=1'b1;
36308: pixelout<=1'b1;
36309: pixelout<=1'b1;
36310: pixelout<=1'b1;
36311: pixelout<=1'b1;
36312: pixelout<=1'b1;
36313: pixelout<=1'b1;
36314: pixelout<=1'b1;
36315: pixelout<=1'b1;
36316: pixelout<=1'b1;
36317: pixelout<=1'b1;
36318: pixelout<=1'b1;
36319: pixelout<=1'b1;
36320: pixelout<=1'b1;
36321: pixelout<=1'b1;
36322: pixelout<=1'b1;
36323: pixelout<=1'b1;
36324: pixelout<=1'b1;
36325: pixelout<=1'b1;
36326: pixelout<=1'b1;
36327: pixelout<=1'b1;
36328: pixelout<=1'b1;
36329: pixelout<=1'b1;
36330: pixelout<=1'b1;
36331: pixelout<=1'b1;
36332: pixelout<=1'b1;
36333: pixelout<=1'b1;
36334: pixelout<=1'b1;
36335: pixelout<=1'b1;
36336: pixelout<=1'b1;
36337: pixelout<=1'b1;
36338: pixelout<=1'b1;
36339: pixelout<=1'b1;
36340: pixelout<=1'b1;
36341: pixelout<=1'b1;
36342: pixelout<=1'b1;
36343: pixelout<=1'b1;
36344: pixelout<=1'b1;
36345: pixelout<=1'b1;
36346: pixelout<=1'b1;
36347: pixelout<=1'b1;
36348: pixelout<=1'b1;
36349: pixelout<=1'b1;
36350: pixelout<=1'b1;
36351: pixelout<=1'b1;
36352: pixelout<=1'b1;
36353: pixelout<=1'b1;
36354: pixelout<=1'b1;
36355: pixelout<=1'b1;
36356: pixelout<=1'b1;
36357: pixelout<=1'b1;
36358: pixelout<=1'b1;
36359: pixelout<=1'b1;
36360: pixelout<=1'b1;
36361: pixelout<=1'b1;
36362: pixelout<=1'b1;
36363: pixelout<=1'b1;
36364: pixelout<=1'b1;
36365: pixelout<=1'b1;
36366: pixelout<=1'b1;
36367: pixelout<=1'b1;
36368: pixelout<=1'b1;
36369: pixelout<=1'b1;
36370: pixelout<=1'b1;
36371: pixelout<=1'b1;
36372: pixelout<=1'b1;
36373: pixelout<=1'b1;
36374: pixelout<=1'b1;
36375: pixelout<=1'b1;
36376: pixelout<=1'b1;
36377: pixelout<=1'b1;
36378: pixelout<=1'b1;
36379: pixelout<=1'b1;
36380: pixelout<=1'b1;
36381: pixelout<=1'b1;
36382: pixelout<=1'b1;
36383: pixelout<=1'b0;
36384: pixelout<=1'b0;
36385: pixelout<=1'b0;
36386: pixelout<=1'b1;
36387: pixelout<=1'b1;
36388: pixelout<=1'b1;
36389: pixelout<=1'b0;
36390: pixelout<=1'b0;
36391: pixelout<=1'b1;
36392: pixelout<=1'b1;
36393: pixelout<=1'b0;
36394: pixelout<=1'b0;
36395: pixelout<=1'b1;
36396: pixelout<=1'b1;
36397: pixelout<=1'b0;
36398: pixelout<=1'b0;
36399: pixelout<=1'b0;
36400: pixelout<=1'b0;
36401: pixelout<=1'b0;
36402: pixelout<=1'b0;
36403: pixelout<=1'b1;
36404: pixelout<=1'b1;
36405: pixelout<=1'b1;
36406: pixelout<=1'b0;
36407: pixelout<=1'b0;
36408: pixelout<=1'b0;
36409: pixelout<=1'b1;
36410: pixelout<=1'b1;
36411: pixelout<=1'b0;
36412: pixelout<=1'b0;
36413: pixelout<=1'b1;
36414: pixelout<=1'b0;
36415: pixelout<=1'b0;
36416: pixelout<=1'b0;
36417: pixelout<=1'b1;
36418: pixelout<=1'b1;
36419: pixelout<=1'b0;
36420: pixelout<=1'b0;
36421: pixelout<=1'b1;
36422: pixelout<=1'b1;
36423: pixelout<=1'b0;
36424: pixelout<=1'b1;
36425: pixelout<=1'b0;
36426: pixelout<=1'b1;
36427: pixelout<=1'b1;
36428: pixelout<=1'b1;
36429: pixelout<=1'b0;
36430: pixelout<=1'b0;
36431: pixelout<=1'b0;
36432: pixelout<=1'b1;
36433: pixelout<=1'b0;
36434: pixelout<=1'b0;
36435: pixelout<=1'b1;
36436: pixelout<=1'b1;
36437: pixelout<=1'b1;
36438: pixelout<=1'b1;
36439: pixelout<=1'b0;
36440: pixelout<=1'b0;
36441: pixelout<=1'b0;
36442: pixelout<=1'b1;
36443: pixelout<=1'b1;
36444: pixelout<=1'b0;
36445: pixelout<=1'b1;
36446: pixelout<=1'b0;
36447: pixelout<=1'b0;
36448: pixelout<=1'b0;
36449: pixelout<=1'b1;
36450: pixelout<=1'b0;
36451: pixelout<=1'b1;
36452: pixelout<=1'b1;
36453: pixelout<=1'b0;
36454: pixelout<=1'b1;
36455: pixelout<=1'b1;
36456: pixelout<=1'b1;
36457: pixelout<=1'b0;
36458: pixelout<=1'b0;
36459: pixelout<=1'b0;
36460: pixelout<=1'b1;
36461: pixelout<=1'b1;
36462: pixelout<=1'b0;
36463: pixelout<=1'b0;
36464: pixelout<=1'b1;
36465: pixelout<=1'b1;
36466: pixelout<=1'b1;
36467: pixelout<=1'b0;
36468: pixelout<=1'b0;
36469: pixelout<=1'b0;
36470: pixelout<=1'b1;
36471: pixelout<=1'b1;
36472: pixelout<=1'b0;
36473: pixelout<=1'b0;
36474: pixelout<=1'b1;
36475: pixelout<=1'b1;
36476: pixelout<=1'b1;
36477: pixelout<=1'b1;
36478: pixelout<=1'b1;
36479: pixelout<=1'b1;
36480: pixelout<=1'b1;
36481: pixelout<=1'b1;
36482: pixelout<=1'b1;
36483: pixelout<=1'b1;
36484: pixelout<=1'b0;
36485: pixelout<=1'b1;
36486: pixelout<=1'b1;
36487: pixelout<=1'b0;
36488: pixelout<=1'b1;
36489: pixelout<=1'b0;
36490: pixelout<=1'b1;
36491: pixelout<=1'b1;
36492: pixelout<=1'b0;
36493: pixelout<=1'b1;
36494: pixelout<=1'b1;
36495: pixelout<=1'b1;
36496: pixelout<=1'b1;
36497: pixelout<=1'b0;
36498: pixelout<=1'b1;
36499: pixelout<=1'b1;
36500: pixelout<=1'b1;
36501: pixelout<=1'b1;
36502: pixelout<=1'b1;
36503: pixelout<=1'b1;
36504: pixelout<=1'b1;
36505: pixelout<=1'b1;
36506: pixelout<=1'b1;
36507: pixelout<=1'b0;
36508: pixelout<=1'b1;
36509: pixelout<=1'b0;
36510: pixelout<=1'b1;
36511: pixelout<=1'b1;
36512: pixelout<=1'b1;
36513: pixelout<=1'b1;
36514: pixelout<=1'b1;
36515: pixelout<=1'b1;
36516: pixelout<=1'b0;
36517: pixelout<=1'b1;
36518: pixelout<=1'b1;
36519: pixelout<=1'b1;
36520: pixelout<=1'b1;
36521: pixelout<=1'b1;
36522: pixelout<=1'b1;
36523: pixelout<=1'b1;
36524: pixelout<=1'b1;
36525: pixelout<=1'b1;
36526: pixelout<=1'b0;
36527: pixelout<=1'b1;
36528: pixelout<=1'b1;
36529: pixelout<=1'b1;
36530: pixelout<=1'b1;
36531: pixelout<=1'b1;
36532: pixelout<=1'b0;
36533: pixelout<=1'b1;
36534: pixelout<=1'b1;
36535: pixelout<=1'b1;
36536: pixelout<=1'b1;
36537: pixelout<=1'b1;
36538: pixelout<=1'b1;
36539: pixelout<=1'b0;
36540: pixelout<=1'b1;
36541: pixelout<=1'b1;
36542: pixelout<=1'b1;
36543: pixelout<=1'b0;
36544: pixelout<=1'b1;
36545: pixelout<=1'b1;
36546: pixelout<=1'b1;
36547: pixelout<=1'b1;
36548: pixelout<=1'b1;
36549: pixelout<=1'b1;
36550: pixelout<=1'b0;
36551: pixelout<=1'b1;
36552: pixelout<=1'b1;
36553: pixelout<=1'b1;
36554: pixelout<=1'b1;
36555: pixelout<=1'b1;
36556: pixelout<=1'b1;
36557: pixelout<=1'b1;
36558: pixelout<=1'b1;
36559: pixelout<=1'b1;
36560: pixelout<=1'b1;
36561: pixelout<=1'b1;
36562: pixelout<=1'b1;
36563: pixelout<=1'b1;
36564: pixelout<=1'b1;
36565: pixelout<=1'b1;
36566: pixelout<=1'b1;
36567: pixelout<=1'b1;
36568: pixelout<=1'b1;
36569: pixelout<=1'b1;
36570: pixelout<=1'b1;
36571: pixelout<=1'b1;
36572: pixelout<=1'b1;
36573: pixelout<=1'b1;
36574: pixelout<=1'b1;
36575: pixelout<=1'b1;
36576: pixelout<=1'b1;
36577: pixelout<=1'b1;
36578: pixelout<=1'b1;
36579: pixelout<=1'b1;
36580: pixelout<=1'b1;
36581: pixelout<=1'b1;
36582: pixelout<=1'b1;
36583: pixelout<=1'b1;
36584: pixelout<=1'b1;
36585: pixelout<=1'b1;
36586: pixelout<=1'b1;
36587: pixelout<=1'b1;
36588: pixelout<=1'b1;
36589: pixelout<=1'b1;
36590: pixelout<=1'b1;
36591: pixelout<=1'b1;
36592: pixelout<=1'b1;
36593: pixelout<=1'b1;
36594: pixelout<=1'b1;
36595: pixelout<=1'b1;
36596: pixelout<=1'b1;
36597: pixelout<=1'b1;
36598: pixelout<=1'b1;
36599: pixelout<=1'b1;
36600: pixelout<=1'b1;
36601: pixelout<=1'b1;
36602: pixelout<=1'b1;
36603: pixelout<=1'b1;
36604: pixelout<=1'b1;
36605: pixelout<=1'b1;
36606: pixelout<=1'b1;
36607: pixelout<=1'b1;
36608: pixelout<=1'b1;
36609: pixelout<=1'b1;
36610: pixelout<=1'b1;
36611: pixelout<=1'b1;
36612: pixelout<=1'b1;
36613: pixelout<=1'b1;
36614: pixelout<=1'b1;
36615: pixelout<=1'b1;
36616: pixelout<=1'b1;
36617: pixelout<=1'b1;
36618: pixelout<=1'b1;
36619: pixelout<=1'b1;
36620: pixelout<=1'b1;
36621: pixelout<=1'b1;
36622: pixelout<=1'b1;
36623: pixelout<=1'b0;
36624: pixelout<=1'b1;
36625: pixelout<=1'b1;
36626: pixelout<=1'b0;
36627: pixelout<=1'b1;
36628: pixelout<=1'b0;
36629: pixelout<=1'b1;
36630: pixelout<=1'b1;
36631: pixelout<=1'b1;
36632: pixelout<=1'b1;
36633: pixelout<=1'b1;
36634: pixelout<=1'b1;
36635: pixelout<=1'b0;
36636: pixelout<=1'b1;
36637: pixelout<=1'b1;
36638: pixelout<=1'b1;
36639: pixelout<=1'b1;
36640: pixelout<=1'b1;
36641: pixelout<=1'b1;
36642: pixelout<=1'b1;
36643: pixelout<=1'b1;
36644: pixelout<=1'b1;
36645: pixelout<=1'b1;
36646: pixelout<=1'b1;
36647: pixelout<=1'b1;
36648: pixelout<=1'b1;
36649: pixelout<=1'b1;
36650: pixelout<=1'b1;
36651: pixelout<=1'b1;
36652: pixelout<=1'b1;
36653: pixelout<=1'b0;
36654: pixelout<=1'b1;
36655: pixelout<=1'b0;
36656: pixelout<=1'b1;
36657: pixelout<=1'b1;
36658: pixelout<=1'b0;
36659: pixelout<=1'b1;
36660: pixelout<=1'b1;
36661: pixelout<=1'b0;
36662: pixelout<=1'b1;
36663: pixelout<=1'b0;
36664: pixelout<=1'b1;
36665: pixelout<=1'b1;
36666: pixelout<=1'b1;
36667: pixelout<=1'b1;
36668: pixelout<=1'b1;
36669: pixelout<=1'b0;
36670: pixelout<=1'b1;
36671: pixelout<=1'b1;
36672: pixelout<=1'b0;
36673: pixelout<=1'b1;
36674: pixelout<=1'b1;
36675: pixelout<=1'b0;
36676: pixelout<=1'b1;
36677: pixelout<=1'b1;
36678: pixelout<=1'b1;
36679: pixelout<=1'b1;
36680: pixelout<=1'b1;
36681: pixelout<=1'b1;
36682: pixelout<=1'b1;
36683: pixelout<=1'b1;
36684: pixelout<=1'b0;
36685: pixelout<=1'b1;
36686: pixelout<=1'b1;
36687: pixelout<=1'b1;
36688: pixelout<=1'b1;
36689: pixelout<=1'b1;
36690: pixelout<=1'b0;
36691: pixelout<=1'b1;
36692: pixelout<=1'b1;
36693: pixelout<=1'b0;
36694: pixelout<=1'b1;
36695: pixelout<=1'b1;
36696: pixelout<=1'b1;
36697: pixelout<=1'b1;
36698: pixelout<=1'b1;
36699: pixelout<=1'b1;
36700: pixelout<=1'b1;
36701: pixelout<=1'b0;
36702: pixelout<=1'b1;
36703: pixelout<=1'b1;
36704: pixelout<=1'b0;
36705: pixelout<=1'b1;
36706: pixelout<=1'b0;
36707: pixelout<=1'b1;
36708: pixelout<=1'b1;
36709: pixelout<=1'b0;
36710: pixelout<=1'b1;
36711: pixelout<=1'b1;
36712: pixelout<=1'b0;
36713: pixelout<=1'b1;
36714: pixelout<=1'b1;
36715: pixelout<=1'b1;
36716: pixelout<=1'b1;
36717: pixelout<=1'b1;
36718: pixelout<=1'b1;
36719: pixelout<=1'b1;
36720: pixelout<=1'b1;
36721: pixelout<=1'b1;
36722: pixelout<=1'b1;
36723: pixelout<=1'b1;
36724: pixelout<=1'b1;
36725: pixelout<=1'b0;
36726: pixelout<=1'b0;
36727: pixelout<=1'b0;
36728: pixelout<=1'b1;
36729: pixelout<=1'b1;
36730: pixelout<=1'b0;
36731: pixelout<=1'b0;
36732: pixelout<=1'b1;
36733: pixelout<=1'b1;
36734: pixelout<=1'b1;
36735: pixelout<=1'b0;
36736: pixelout<=1'b0;
36737: pixelout<=1'b1;
36738: pixelout<=1'b1;
36739: pixelout<=1'b0;
36740: pixelout<=1'b0;
36741: pixelout<=1'b0;
36742: pixelout<=1'b1;
36743: pixelout<=1'b1;
36744: pixelout<=1'b1;
36745: pixelout<=1'b1;
36746: pixelout<=1'b1;
36747: pixelout<=1'b1;
36748: pixelout<=1'b0;
36749: pixelout<=1'b1;
36750: pixelout<=1'b0;
36751: pixelout<=1'b1;
36752: pixelout<=1'b1;
36753: pixelout<=1'b0;
36754: pixelout<=1'b0;
36755: pixelout<=1'b1;
36756: pixelout<=1'b0;
36757: pixelout<=1'b1;
36758: pixelout<=1'b1;
36759: pixelout<=1'b1;
36760: pixelout<=1'b1;
36761: pixelout<=1'b1;
36762: pixelout<=1'b1;
36763: pixelout<=1'b1;
36764: pixelout<=1'b1;
36765: pixelout<=1'b1;
36766: pixelout<=1'b0;
36767: pixelout<=1'b1;
36768: pixelout<=1'b1;
36769: pixelout<=1'b1;
36770: pixelout<=1'b0;
36771: pixelout<=1'b0;
36772: pixelout<=1'b1;
36773: pixelout<=1'b1;
36774: pixelout<=1'b0;
36775: pixelout<=1'b0;
36776: pixelout<=1'b0;
36777: pixelout<=1'b1;
36778: pixelout<=1'b1;
36779: pixelout<=1'b0;
36780: pixelout<=1'b1;
36781: pixelout<=1'b1;
36782: pixelout<=1'b1;
36783: pixelout<=1'b1;
36784: pixelout<=1'b1;
36785: pixelout<=1'b1;
36786: pixelout<=1'b1;
36787: pixelout<=1'b1;
36788: pixelout<=1'b1;
36789: pixelout<=1'b1;
36790: pixelout<=1'b1;
36791: pixelout<=1'b1;
36792: pixelout<=1'b1;
36793: pixelout<=1'b1;
36794: pixelout<=1'b1;
36795: pixelout<=1'b1;
36796: pixelout<=1'b1;
36797: pixelout<=1'b1;
36798: pixelout<=1'b1;
36799: pixelout<=1'b1;
36800: pixelout<=1'b1;
36801: pixelout<=1'b1;
36802: pixelout<=1'b1;
36803: pixelout<=1'b1;
36804: pixelout<=1'b1;
36805: pixelout<=1'b1;
36806: pixelout<=1'b1;
36807: pixelout<=1'b1;
36808: pixelout<=1'b1;
36809: pixelout<=1'b1;
36810: pixelout<=1'b1;
36811: pixelout<=1'b1;
36812: pixelout<=1'b1;
36813: pixelout<=1'b1;
36814: pixelout<=1'b1;
36815: pixelout<=1'b1;
36816: pixelout<=1'b1;
36817: pixelout<=1'b1;
36818: pixelout<=1'b1;
36819: pixelout<=1'b1;
36820: pixelout<=1'b1;
36821: pixelout<=1'b1;
36822: pixelout<=1'b1;
36823: pixelout<=1'b1;
36824: pixelout<=1'b1;
36825: pixelout<=1'b1;
36826: pixelout<=1'b1;
36827: pixelout<=1'b1;
36828: pixelout<=1'b1;
36829: pixelout<=1'b1;
36830: pixelout<=1'b1;
36831: pixelout<=1'b1;
36832: pixelout<=1'b1;
36833: pixelout<=1'b1;
36834: pixelout<=1'b1;
36835: pixelout<=1'b1;
36836: pixelout<=1'b1;
36837: pixelout<=1'b1;
36838: pixelout<=1'b1;
36839: pixelout<=1'b1;
36840: pixelout<=1'b1;
36841: pixelout<=1'b1;
36842: pixelout<=1'b1;
36843: pixelout<=1'b1;
36844: pixelout<=1'b1;
36845: pixelout<=1'b1;
36846: pixelout<=1'b1;
36847: pixelout<=1'b1;
36848: pixelout<=1'b1;
36849: pixelout<=1'b1;
36850: pixelout<=1'b1;
36851: pixelout<=1'b1;
36852: pixelout<=1'b1;
36853: pixelout<=1'b1;
36854: pixelout<=1'b1;
36855: pixelout<=1'b1;
36856: pixelout<=1'b1;
36857: pixelout<=1'b1;
36858: pixelout<=1'b1;
36859: pixelout<=1'b1;
36860: pixelout<=1'b1;
36861: pixelout<=1'b1;
36862: pixelout<=1'b1;
36863: pixelout<=1'b0;
36864: pixelout<=1'b1;
36865: pixelout<=1'b1;
36866: pixelout<=1'b0;
36867: pixelout<=1'b1;
36868: pixelout<=1'b1;
36869: pixelout<=1'b1;
36870: pixelout<=1'b1;
36871: pixelout<=1'b1;
36872: pixelout<=1'b0;
36873: pixelout<=1'b1;
36874: pixelout<=1'b1;
36875: pixelout<=1'b1;
36876: pixelout<=1'b1;
36877: pixelout<=1'b1;
36878: pixelout<=1'b1;
36879: pixelout<=1'b1;
36880: pixelout<=1'b1;
36881: pixelout<=1'b1;
36882: pixelout<=1'b1;
36883: pixelout<=1'b1;
36884: pixelout<=1'b1;
36885: pixelout<=1'b1;
36886: pixelout<=1'b1;
36887: pixelout<=1'b1;
36888: pixelout<=1'b1;
36889: pixelout<=1'b1;
36890: pixelout<=1'b1;
36891: pixelout<=1'b1;
36892: pixelout<=1'b1;
36893: pixelout<=1'b0;
36894: pixelout<=1'b1;
36895: pixelout<=1'b0;
36896: pixelout<=1'b1;
36897: pixelout<=1'b1;
36898: pixelout<=1'b0;
36899: pixelout<=1'b1;
36900: pixelout<=1'b1;
36901: pixelout<=1'b1;
36902: pixelout<=1'b1;
36903: pixelout<=1'b0;
36904: pixelout<=1'b1;
36905: pixelout<=1'b1;
36906: pixelout<=1'b1;
36907: pixelout<=1'b1;
36908: pixelout<=1'b1;
36909: pixelout<=1'b0;
36910: pixelout<=1'b1;
36911: pixelout<=1'b1;
36912: pixelout<=1'b0;
36913: pixelout<=1'b1;
36914: pixelout<=1'b1;
36915: pixelout<=1'b0;
36916: pixelout<=1'b1;
36917: pixelout<=1'b1;
36918: pixelout<=1'b1;
36919: pixelout<=1'b1;
36920: pixelout<=1'b1;
36921: pixelout<=1'b1;
36922: pixelout<=1'b1;
36923: pixelout<=1'b1;
36924: pixelout<=1'b0;
36925: pixelout<=1'b1;
36926: pixelout<=1'b1;
36927: pixelout<=1'b1;
36928: pixelout<=1'b0;
36929: pixelout<=1'b1;
36930: pixelout<=1'b0;
36931: pixelout<=1'b1;
36932: pixelout<=1'b1;
36933: pixelout<=1'b0;
36934: pixelout<=1'b1;
36935: pixelout<=1'b1;
36936: pixelout<=1'b1;
36937: pixelout<=1'b1;
36938: pixelout<=1'b1;
36939: pixelout<=1'b0;
36940: pixelout<=1'b1;
36941: pixelout<=1'b0;
36942: pixelout<=1'b1;
36943: pixelout<=1'b1;
36944: pixelout<=1'b0;
36945: pixelout<=1'b1;
36946: pixelout<=1'b0;
36947: pixelout<=1'b1;
36948: pixelout<=1'b1;
36949: pixelout<=1'b0;
36950: pixelout<=1'b1;
36951: pixelout<=1'b1;
36952: pixelout<=1'b0;
36953: pixelout<=1'b1;
36954: pixelout<=1'b1;
36955: pixelout<=1'b1;
36956: pixelout<=1'b1;
36957: pixelout<=1'b1;
36958: pixelout<=1'b1;
36959: pixelout<=1'b1;
36960: pixelout<=1'b1;
36961: pixelout<=1'b1;
36962: pixelout<=1'b1;
36963: pixelout<=1'b1;
36964: pixelout<=1'b1;
36965: pixelout<=1'b1;
36966: pixelout<=1'b1;
36967: pixelout<=1'b0;
36968: pixelout<=1'b1;
36969: pixelout<=1'b1;
36970: pixelout<=1'b1;
36971: pixelout<=1'b1;
36972: pixelout<=1'b1;
36973: pixelout<=1'b1;
36974: pixelout<=1'b1;
36975: pixelout<=1'b1;
36976: pixelout<=1'b1;
36977: pixelout<=1'b1;
36978: pixelout<=1'b1;
36979: pixelout<=1'b1;
36980: pixelout<=1'b1;
36981: pixelout<=1'b1;
36982: pixelout<=1'b1;
36983: pixelout<=1'b1;
36984: pixelout<=1'b1;
36985: pixelout<=1'b1;
36986: pixelout<=1'b1;
36987: pixelout<=1'b1;
36988: pixelout<=1'b1;
36989: pixelout<=1'b1;
36990: pixelout<=1'b1;
36991: pixelout<=1'b1;
36992: pixelout<=1'b1;
36993: pixelout<=1'b1;
36994: pixelout<=1'b1;
36995: pixelout<=1'b1;
36996: pixelout<=1'b1;
36997: pixelout<=1'b1;
36998: pixelout<=1'b1;
36999: pixelout<=1'b1;
37000: pixelout<=1'b1;
37001: pixelout<=1'b1;
37002: pixelout<=1'b1;
37003: pixelout<=1'b1;
37004: pixelout<=1'b1;
37005: pixelout<=1'b1;
37006: pixelout<=1'b1;
37007: pixelout<=1'b1;
37008: pixelout<=1'b1;
37009: pixelout<=1'b1;
37010: pixelout<=1'b1;
37011: pixelout<=1'b1;
37012: pixelout<=1'b1;
37013: pixelout<=1'b1;
37014: pixelout<=1'b1;
37015: pixelout<=1'b1;
37016: pixelout<=1'b1;
37017: pixelout<=1'b1;
37018: pixelout<=1'b1;
37019: pixelout<=1'b1;
37020: pixelout<=1'b1;
37021: pixelout<=1'b1;
37022: pixelout<=1'b1;
37023: pixelout<=1'b1;
37024: pixelout<=1'b1;
37025: pixelout<=1'b1;
37026: pixelout<=1'b1;
37027: pixelout<=1'b1;
37028: pixelout<=1'b1;
37029: pixelout<=1'b1;
37030: pixelout<=1'b1;
37031: pixelout<=1'b1;
37032: pixelout<=1'b1;
37033: pixelout<=1'b1;
37034: pixelout<=1'b1;
37035: pixelout<=1'b1;
37036: pixelout<=1'b1;
37037: pixelout<=1'b1;
37038: pixelout<=1'b1;
37039: pixelout<=1'b1;
37040: pixelout<=1'b1;
37041: pixelout<=1'b1;
37042: pixelout<=1'b1;
37043: pixelout<=1'b1;
37044: pixelout<=1'b1;
37045: pixelout<=1'b1;
37046: pixelout<=1'b1;
37047: pixelout<=1'b1;
37048: pixelout<=1'b1;
37049: pixelout<=1'b1;
37050: pixelout<=1'b1;
37051: pixelout<=1'b1;
37052: pixelout<=1'b1;
37053: pixelout<=1'b1;
37054: pixelout<=1'b1;
37055: pixelout<=1'b1;
37056: pixelout<=1'b1;
37057: pixelout<=1'b1;
37058: pixelout<=1'b1;
37059: pixelout<=1'b1;
37060: pixelout<=1'b1;
37061: pixelout<=1'b1;
37062: pixelout<=1'b1;
37063: pixelout<=1'b1;
37064: pixelout<=1'b1;
37065: pixelout<=1'b1;
37066: pixelout<=1'b1;
37067: pixelout<=1'b1;
37068: pixelout<=1'b1;
37069: pixelout<=1'b1;
37070: pixelout<=1'b1;
37071: pixelout<=1'b1;
37072: pixelout<=1'b1;
37073: pixelout<=1'b1;
37074: pixelout<=1'b1;
37075: pixelout<=1'b1;
37076: pixelout<=1'b1;
37077: pixelout<=1'b1;
37078: pixelout<=1'b1;
37079: pixelout<=1'b1;
37080: pixelout<=1'b1;
37081: pixelout<=1'b1;
37082: pixelout<=1'b1;
37083: pixelout<=1'b1;
37084: pixelout<=1'b1;
37085: pixelout<=1'b1;
37086: pixelout<=1'b1;
37087: pixelout<=1'b1;
37088: pixelout<=1'b1;
37089: pixelout<=1'b1;
37090: pixelout<=1'b1;
37091: pixelout<=1'b1;
37092: pixelout<=1'b1;
37093: pixelout<=1'b1;
37094: pixelout<=1'b1;
37095: pixelout<=1'b1;
37096: pixelout<=1'b1;
37097: pixelout<=1'b1;
37098: pixelout<=1'b1;
37099: pixelout<=1'b1;
37100: pixelout<=1'b1;
37101: pixelout<=1'b1;
37102: pixelout<=1'b1;
37103: pixelout<=1'b0;
37104: pixelout<=1'b0;
37105: pixelout<=1'b0;
37106: pixelout<=1'b1;
37107: pixelout<=1'b1;
37108: pixelout<=1'b1;
37109: pixelout<=1'b1;
37110: pixelout<=1'b1;
37111: pixelout<=1'b1;
37112: pixelout<=1'b1;
37113: pixelout<=1'b0;
37114: pixelout<=1'b0;
37115: pixelout<=1'b1;
37116: pixelout<=1'b1;
37117: pixelout<=1'b0;
37118: pixelout<=1'b0;
37119: pixelout<=1'b0;
37120: pixelout<=1'b1;
37121: pixelout<=1'b0;
37122: pixelout<=1'b0;
37123: pixelout<=1'b1;
37124: pixelout<=1'b1;
37125: pixelout<=1'b1;
37126: pixelout<=1'b0;
37127: pixelout<=1'b0;
37128: pixelout<=1'b0;
37129: pixelout<=1'b1;
37130: pixelout<=1'b1;
37131: pixelout<=1'b1;
37132: pixelout<=1'b1;
37133: pixelout<=1'b0;
37134: pixelout<=1'b1;
37135: pixelout<=1'b0;
37136: pixelout<=1'b0;
37137: pixelout<=1'b1;
37138: pixelout<=1'b1;
37139: pixelout<=1'b0;
37140: pixelout<=1'b0;
37141: pixelout<=1'b0;
37142: pixelout<=1'b1;
37143: pixelout<=1'b0;
37144: pixelout<=1'b1;
37145: pixelout<=1'b1;
37146: pixelout<=1'b1;
37147: pixelout<=1'b1;
37148: pixelout<=1'b1;
37149: pixelout<=1'b0;
37150: pixelout<=1'b0;
37151: pixelout<=1'b1;
37152: pixelout<=1'b1;
37153: pixelout<=1'b0;
37154: pixelout<=1'b0;
37155: pixelout<=1'b1;
37156: pixelout<=1'b1;
37157: pixelout<=1'b1;
37158: pixelout<=1'b1;
37159: pixelout<=1'b0;
37160: pixelout<=1'b0;
37161: pixelout<=1'b0;
37162: pixelout<=1'b1;
37163: pixelout<=1'b1;
37164: pixelout<=1'b0;
37165: pixelout<=1'b1;
37166: pixelout<=1'b0;
37167: pixelout<=1'b0;
37168: pixelout<=1'b1;
37169: pixelout<=1'b1;
37170: pixelout<=1'b1;
37171: pixelout<=1'b0;
37172: pixelout<=1'b0;
37173: pixelout<=1'b0;
37174: pixelout<=1'b1;
37175: pixelout<=1'b1;
37176: pixelout<=1'b1;
37177: pixelout<=1'b0;
37178: pixelout<=1'b0;
37179: pixelout<=1'b1;
37180: pixelout<=1'b1;
37181: pixelout<=1'b1;
37182: pixelout<=1'b0;
37183: pixelout<=1'b0;
37184: pixelout<=1'b0;
37185: pixelout<=1'b1;
37186: pixelout<=1'b1;
37187: pixelout<=1'b0;
37188: pixelout<=1'b1;
37189: pixelout<=1'b0;
37190: pixelout<=1'b1;
37191: pixelout<=1'b1;
37192: pixelout<=1'b0;
37193: pixelout<=1'b1;
37194: pixelout<=1'b1;
37195: pixelout<=1'b1;
37196: pixelout<=1'b1;
37197: pixelout<=1'b1;
37198: pixelout<=1'b1;
37199: pixelout<=1'b1;
37200: pixelout<=1'b1;
37201: pixelout<=1'b1;
37202: pixelout<=1'b1;
37203: pixelout<=1'b1;
37204: pixelout<=1'b1;
37205: pixelout<=1'b1;
37206: pixelout<=1'b1;
37207: pixelout<=1'b1;
37208: pixelout<=1'b1;
37209: pixelout<=1'b1;
37210: pixelout<=1'b1;
37211: pixelout<=1'b1;
37212: pixelout<=1'b1;
37213: pixelout<=1'b1;
37214: pixelout<=1'b1;
37215: pixelout<=1'b1;
37216: pixelout<=1'b1;
37217: pixelout<=1'b1;
37218: pixelout<=1'b1;
37219: pixelout<=1'b1;
37220: pixelout<=1'b1;
37221: pixelout<=1'b1;
37222: pixelout<=1'b1;
37223: pixelout<=1'b1;
37224: pixelout<=1'b1;
37225: pixelout<=1'b1;
37226: pixelout<=1'b1;
37227: pixelout<=1'b1;
37228: pixelout<=1'b1;
37229: pixelout<=1'b1;
37230: pixelout<=1'b1;
37231: pixelout<=1'b1;
37232: pixelout<=1'b1;
37233: pixelout<=1'b1;
37234: pixelout<=1'b1;
37235: pixelout<=1'b1;
37236: pixelout<=1'b1;
37237: pixelout<=1'b1;
37238: pixelout<=1'b1;
37239: pixelout<=1'b1;
37240: pixelout<=1'b1;
37241: pixelout<=1'b1;
37242: pixelout<=1'b1;
37243: pixelout<=1'b1;
37244: pixelout<=1'b1;
37245: pixelout<=1'b1;
37246: pixelout<=1'b1;
37247: pixelout<=1'b1;
37248: pixelout<=1'b1;
37249: pixelout<=1'b1;
37250: pixelout<=1'b1;
37251: pixelout<=1'b1;
37252: pixelout<=1'b1;
37253: pixelout<=1'b1;
37254: pixelout<=1'b1;
37255: pixelout<=1'b1;
37256: pixelout<=1'b1;
37257: pixelout<=1'b1;
37258: pixelout<=1'b1;
37259: pixelout<=1'b1;
37260: pixelout<=1'b1;
37261: pixelout<=1'b1;
37262: pixelout<=1'b1;
37263: pixelout<=1'b1;
37264: pixelout<=1'b1;
37265: pixelout<=1'b1;
37266: pixelout<=1'b1;
37267: pixelout<=1'b1;
37268: pixelout<=1'b1;
37269: pixelout<=1'b1;
37270: pixelout<=1'b1;
37271: pixelout<=1'b1;
37272: pixelout<=1'b1;
37273: pixelout<=1'b1;
37274: pixelout<=1'b1;
37275: pixelout<=1'b1;
37276: pixelout<=1'b1;
37277: pixelout<=1'b1;
37278: pixelout<=1'b1;
37279: pixelout<=1'b1;
37280: pixelout<=1'b1;
37281: pixelout<=1'b1;
37282: pixelout<=1'b1;
37283: pixelout<=1'b1;
37284: pixelout<=1'b1;
37285: pixelout<=1'b1;
37286: pixelout<=1'b1;
37287: pixelout<=1'b1;
37288: pixelout<=1'b1;
37289: pixelout<=1'b1;
37290: pixelout<=1'b1;
37291: pixelout<=1'b1;
37292: pixelout<=1'b1;
37293: pixelout<=1'b1;
37294: pixelout<=1'b1;
37295: pixelout<=1'b1;
37296: pixelout<=1'b1;
37297: pixelout<=1'b1;
37298: pixelout<=1'b1;
37299: pixelout<=1'b1;
37300: pixelout<=1'b1;
37301: pixelout<=1'b1;
37302: pixelout<=1'b1;
37303: pixelout<=1'b1;
37304: pixelout<=1'b1;
37305: pixelout<=1'b1;
37306: pixelout<=1'b1;
37307: pixelout<=1'b1;
37308: pixelout<=1'b1;
37309: pixelout<=1'b1;
37310: pixelout<=1'b1;
37311: pixelout<=1'b1;
37312: pixelout<=1'b1;
37313: pixelout<=1'b1;
37314: pixelout<=1'b1;
37315: pixelout<=1'b1;
37316: pixelout<=1'b1;
37317: pixelout<=1'b1;
37318: pixelout<=1'b1;
37319: pixelout<=1'b1;
37320: pixelout<=1'b1;
37321: pixelout<=1'b1;
37322: pixelout<=1'b1;
37323: pixelout<=1'b1;
37324: pixelout<=1'b1;
37325: pixelout<=1'b1;
37326: pixelout<=1'b1;
37327: pixelout<=1'b1;
37328: pixelout<=1'b1;
37329: pixelout<=1'b1;
37330: pixelout<=1'b1;
37331: pixelout<=1'b1;
37332: pixelout<=1'b1;
37333: pixelout<=1'b1;
37334: pixelout<=1'b1;
37335: pixelout<=1'b1;
37336: pixelout<=1'b1;
37337: pixelout<=1'b1;
37338: pixelout<=1'b1;
37339: pixelout<=1'b1;
37340: pixelout<=1'b1;
37341: pixelout<=1'b1;
37342: pixelout<=1'b1;
37343: pixelout<=1'b0;
37344: pixelout<=1'b1;
37345: pixelout<=1'b1;
37346: pixelout<=1'b1;
37347: pixelout<=1'b1;
37348: pixelout<=1'b1;
37349: pixelout<=1'b1;
37350: pixelout<=1'b1;
37351: pixelout<=1'b1;
37352: pixelout<=1'b1;
37353: pixelout<=1'b1;
37354: pixelout<=1'b1;
37355: pixelout<=1'b1;
37356: pixelout<=1'b1;
37357: pixelout<=1'b1;
37358: pixelout<=1'b1;
37359: pixelout<=1'b1;
37360: pixelout<=1'b1;
37361: pixelout<=1'b1;
37362: pixelout<=1'b1;
37363: pixelout<=1'b1;
37364: pixelout<=1'b1;
37365: pixelout<=1'b1;
37366: pixelout<=1'b1;
37367: pixelout<=1'b1;
37368: pixelout<=1'b1;
37369: pixelout<=1'b1;
37370: pixelout<=1'b1;
37371: pixelout<=1'b1;
37372: pixelout<=1'b1;
37373: pixelout<=1'b1;
37374: pixelout<=1'b1;
37375: pixelout<=1'b1;
37376: pixelout<=1'b1;
37377: pixelout<=1'b1;
37378: pixelout<=1'b1;
37379: pixelout<=1'b1;
37380: pixelout<=1'b1;
37381: pixelout<=1'b1;
37382: pixelout<=1'b1;
37383: pixelout<=1'b1;
37384: pixelout<=1'b1;
37385: pixelout<=1'b1;
37386: pixelout<=1'b1;
37387: pixelout<=1'b1;
37388: pixelout<=1'b1;
37389: pixelout<=1'b1;
37390: pixelout<=1'b1;
37391: pixelout<=1'b1;
37392: pixelout<=1'b1;
37393: pixelout<=1'b1;
37394: pixelout<=1'b1;
37395: pixelout<=1'b1;
37396: pixelout<=1'b1;
37397: pixelout<=1'b1;
37398: pixelout<=1'b1;
37399: pixelout<=1'b1;
37400: pixelout<=1'b1;
37401: pixelout<=1'b1;
37402: pixelout<=1'b1;
37403: pixelout<=1'b1;
37404: pixelout<=1'b1;
37405: pixelout<=1'b1;
37406: pixelout<=1'b1;
37407: pixelout<=1'b1;
37408: pixelout<=1'b1;
37409: pixelout<=1'b1;
37410: pixelout<=1'b1;
37411: pixelout<=1'b1;
37412: pixelout<=1'b1;
37413: pixelout<=1'b0;
37414: pixelout<=1'b1;
37415: pixelout<=1'b1;
37416: pixelout<=1'b1;
37417: pixelout<=1'b1;
37418: pixelout<=1'b1;
37419: pixelout<=1'b1;
37420: pixelout<=1'b1;
37421: pixelout<=1'b1;
37422: pixelout<=1'b1;
37423: pixelout<=1'b1;
37424: pixelout<=1'b0;
37425: pixelout<=1'b1;
37426: pixelout<=1'b1;
37427: pixelout<=1'b1;
37428: pixelout<=1'b1;
37429: pixelout<=1'b1;
37430: pixelout<=1'b1;
37431: pixelout<=1'b1;
37432: pixelout<=1'b1;
37433: pixelout<=1'b1;
37434: pixelout<=1'b1;
37435: pixelout<=1'b1;
37436: pixelout<=1'b1;
37437: pixelout<=1'b1;
37438: pixelout<=1'b1;
37439: pixelout<=1'b1;
37440: pixelout<=1'b1;
37441: pixelout<=1'b1;
37442: pixelout<=1'b1;
37443: pixelout<=1'b1;
37444: pixelout<=1'b1;
37445: pixelout<=1'b1;
37446: pixelout<=1'b1;
37447: pixelout<=1'b1;
37448: pixelout<=1'b1;
37449: pixelout<=1'b1;
37450: pixelout<=1'b1;
37451: pixelout<=1'b1;
37452: pixelout<=1'b1;
37453: pixelout<=1'b1;
37454: pixelout<=1'b1;
37455: pixelout<=1'b1;
37456: pixelout<=1'b1;
37457: pixelout<=1'b1;
37458: pixelout<=1'b1;
37459: pixelout<=1'b1;
37460: pixelout<=1'b1;
37461: pixelout<=1'b1;
37462: pixelout<=1'b1;
37463: pixelout<=1'b1;
37464: pixelout<=1'b1;
37465: pixelout<=1'b1;
37466: pixelout<=1'b1;
37467: pixelout<=1'b1;
37468: pixelout<=1'b1;
37469: pixelout<=1'b1;
37470: pixelout<=1'b1;
37471: pixelout<=1'b1;
37472: pixelout<=1'b1;
37473: pixelout<=1'b1;
37474: pixelout<=1'b1;
37475: pixelout<=1'b1;
37476: pixelout<=1'b1;
37477: pixelout<=1'b1;
37478: pixelout<=1'b1;
37479: pixelout<=1'b1;
37480: pixelout<=1'b1;
37481: pixelout<=1'b1;
37482: pixelout<=1'b1;
37483: pixelout<=1'b1;
37484: pixelout<=1'b1;
37485: pixelout<=1'b1;
37486: pixelout<=1'b1;
37487: pixelout<=1'b1;
37488: pixelout<=1'b1;
37489: pixelout<=1'b1;
37490: pixelout<=1'b1;
37491: pixelout<=1'b1;
37492: pixelout<=1'b1;
37493: pixelout<=1'b1;
37494: pixelout<=1'b1;
37495: pixelout<=1'b1;
37496: pixelout<=1'b1;
37497: pixelout<=1'b1;
37498: pixelout<=1'b1;
37499: pixelout<=1'b1;
37500: pixelout<=1'b1;
37501: pixelout<=1'b1;
37502: pixelout<=1'b1;
37503: pixelout<=1'b1;
37504: pixelout<=1'b1;
37505: pixelout<=1'b1;
37506: pixelout<=1'b1;
37507: pixelout<=1'b1;
37508: pixelout<=1'b1;
37509: pixelout<=1'b1;
37510: pixelout<=1'b1;
37511: pixelout<=1'b1;
37512: pixelout<=1'b1;
37513: pixelout<=1'b1;
37514: pixelout<=1'b1;
37515: pixelout<=1'b1;
37516: pixelout<=1'b1;
37517: pixelout<=1'b1;
37518: pixelout<=1'b1;
37519: pixelout<=1'b1;
37520: pixelout<=1'b1;
37521: pixelout<=1'b1;
37522: pixelout<=1'b1;
37523: pixelout<=1'b1;
37524: pixelout<=1'b1;
37525: pixelout<=1'b1;
37526: pixelout<=1'b1;
37527: pixelout<=1'b1;
37528: pixelout<=1'b1;
37529: pixelout<=1'b1;
37530: pixelout<=1'b1;
37531: pixelout<=1'b1;
37532: pixelout<=1'b1;
37533: pixelout<=1'b1;
37534: pixelout<=1'b1;
37535: pixelout<=1'b1;
37536: pixelout<=1'b1;
37537: pixelout<=1'b1;
37538: pixelout<=1'b1;
37539: pixelout<=1'b1;
37540: pixelout<=1'b1;
37541: pixelout<=1'b1;
37542: pixelout<=1'b1;
37543: pixelout<=1'b1;
37544: pixelout<=1'b1;
37545: pixelout<=1'b1;
37546: pixelout<=1'b1;
37547: pixelout<=1'b1;
37548: pixelout<=1'b1;
37549: pixelout<=1'b1;
37550: pixelout<=1'b1;
37551: pixelout<=1'b1;
37552: pixelout<=1'b1;
37553: pixelout<=1'b1;
37554: pixelout<=1'b1;
37555: pixelout<=1'b1;
37556: pixelout<=1'b1;
37557: pixelout<=1'b1;
37558: pixelout<=1'b1;
37559: pixelout<=1'b1;
37560: pixelout<=1'b1;
37561: pixelout<=1'b1;
37562: pixelout<=1'b1;
37563: pixelout<=1'b1;
37564: pixelout<=1'b1;
37565: pixelout<=1'b1;
37566: pixelout<=1'b1;
37567: pixelout<=1'b1;
37568: pixelout<=1'b1;
37569: pixelout<=1'b1;
37570: pixelout<=1'b1;
37571: pixelout<=1'b1;
37572: pixelout<=1'b1;
37573: pixelout<=1'b1;
37574: pixelout<=1'b1;
37575: pixelout<=1'b1;
37576: pixelout<=1'b1;
37577: pixelout<=1'b1;
37578: pixelout<=1'b1;
37579: pixelout<=1'b1;
37580: pixelout<=1'b1;
37581: pixelout<=1'b1;
37582: pixelout<=1'b1;
37583: pixelout<=1'b1;
37584: pixelout<=1'b1;
37585: pixelout<=1'b1;
37586: pixelout<=1'b1;
37587: pixelout<=1'b1;
37588: pixelout<=1'b1;
37589: pixelout<=1'b1;
37590: pixelout<=1'b1;
37591: pixelout<=1'b1;
37592: pixelout<=1'b1;
37593: pixelout<=1'b1;
37594: pixelout<=1'b1;
37595: pixelout<=1'b1;
37596: pixelout<=1'b1;
37597: pixelout<=1'b1;
37598: pixelout<=1'b1;
37599: pixelout<=1'b1;
37600: pixelout<=1'b1;
37601: pixelout<=1'b1;
37602: pixelout<=1'b1;
37603: pixelout<=1'b1;
37604: pixelout<=1'b1;
37605: pixelout<=1'b1;
37606: pixelout<=1'b1;
37607: pixelout<=1'b1;
37608: pixelout<=1'b1;
37609: pixelout<=1'b1;
37610: pixelout<=1'b1;
37611: pixelout<=1'b1;
37612: pixelout<=1'b1;
37613: pixelout<=1'b1;
37614: pixelout<=1'b1;
37615: pixelout<=1'b1;
37616: pixelout<=1'b1;
37617: pixelout<=1'b1;
37618: pixelout<=1'b1;
37619: pixelout<=1'b1;
37620: pixelout<=1'b1;
37621: pixelout<=1'b1;
37622: pixelout<=1'b1;
37623: pixelout<=1'b1;
37624: pixelout<=1'b1;
37625: pixelout<=1'b1;
37626: pixelout<=1'b1;
37627: pixelout<=1'b1;
37628: pixelout<=1'b1;
37629: pixelout<=1'b1;
37630: pixelout<=1'b1;
37631: pixelout<=1'b1;
37632: pixelout<=1'b1;
37633: pixelout<=1'b1;
37634: pixelout<=1'b1;
37635: pixelout<=1'b1;
37636: pixelout<=1'b1;
37637: pixelout<=1'b1;
37638: pixelout<=1'b1;
37639: pixelout<=1'b1;
37640: pixelout<=1'b1;
37641: pixelout<=1'b1;
37642: pixelout<=1'b1;
37643: pixelout<=1'b1;
37644: pixelout<=1'b1;
37645: pixelout<=1'b1;
37646: pixelout<=1'b1;
37647: pixelout<=1'b1;
37648: pixelout<=1'b1;
37649: pixelout<=1'b1;
37650: pixelout<=1'b1;
37651: pixelout<=1'b1;
37652: pixelout<=1'b1;
37653: pixelout<=1'b1;
37654: pixelout<=1'b1;
37655: pixelout<=1'b1;
37656: pixelout<=1'b1;
37657: pixelout<=1'b1;
37658: pixelout<=1'b1;
37659: pixelout<=1'b1;
37660: pixelout<=1'b1;
37661: pixelout<=1'b1;
37662: pixelout<=1'b1;
37663: pixelout<=1'b1;
37664: pixelout<=1'b1;
37665: pixelout<=1'b1;
37666: pixelout<=1'b1;
37667: pixelout<=1'b1;
37668: pixelout<=1'b1;
37669: pixelout<=1'b1;
37670: pixelout<=1'b1;
37671: pixelout<=1'b1;
37672: pixelout<=1'b1;
37673: pixelout<=1'b1;
37674: pixelout<=1'b1;
37675: pixelout<=1'b1;
37676: pixelout<=1'b1;
37677: pixelout<=1'b1;
37678: pixelout<=1'b1;
37679: pixelout<=1'b1;
37680: pixelout<=1'b1;
37681: pixelout<=1'b1;
37682: pixelout<=1'b1;
37683: pixelout<=1'b1;
37684: pixelout<=1'b1;
37685: pixelout<=1'b1;
37686: pixelout<=1'b1;
37687: pixelout<=1'b1;
37688: pixelout<=1'b1;
37689: pixelout<=1'b1;
37690: pixelout<=1'b1;
37691: pixelout<=1'b1;
37692: pixelout<=1'b1;
37693: pixelout<=1'b1;
37694: pixelout<=1'b1;
37695: pixelout<=1'b1;
37696: pixelout<=1'b1;
37697: pixelout<=1'b1;
37698: pixelout<=1'b1;
37699: pixelout<=1'b1;
37700: pixelout<=1'b1;
37701: pixelout<=1'b1;
37702: pixelout<=1'b1;
37703: pixelout<=1'b1;
37704: pixelout<=1'b1;
37705: pixelout<=1'b1;
37706: pixelout<=1'b1;
37707: pixelout<=1'b1;
37708: pixelout<=1'b1;
37709: pixelout<=1'b1;
37710: pixelout<=1'b1;
37711: pixelout<=1'b1;
37712: pixelout<=1'b1;
37713: pixelout<=1'b1;
37714: pixelout<=1'b1;
37715: pixelout<=1'b1;
37716: pixelout<=1'b1;
37717: pixelout<=1'b1;
37718: pixelout<=1'b1;
37719: pixelout<=1'b1;
37720: pixelout<=1'b1;
37721: pixelout<=1'b1;
37722: pixelout<=1'b1;
37723: pixelout<=1'b1;
37724: pixelout<=1'b1;
37725: pixelout<=1'b1;
37726: pixelout<=1'b1;
37727: pixelout<=1'b1;
37728: pixelout<=1'b1;
37729: pixelout<=1'b1;
37730: pixelout<=1'b1;
37731: pixelout<=1'b1;
37732: pixelout<=1'b1;
37733: pixelout<=1'b1;
37734: pixelout<=1'b1;
37735: pixelout<=1'b1;
37736: pixelout<=1'b1;
37737: pixelout<=1'b1;
37738: pixelout<=1'b1;
37739: pixelout<=1'b1;
37740: pixelout<=1'b1;
37741: pixelout<=1'b1;
37742: pixelout<=1'b1;
37743: pixelout<=1'b1;
37744: pixelout<=1'b1;
37745: pixelout<=1'b1;
37746: pixelout<=1'b1;
37747: pixelout<=1'b1;
37748: pixelout<=1'b1;
37749: pixelout<=1'b1;
37750: pixelout<=1'b1;
37751: pixelout<=1'b1;
37752: pixelout<=1'b1;
37753: pixelout<=1'b1;
37754: pixelout<=1'b1;
37755: pixelout<=1'b1;
37756: pixelout<=1'b1;
37757: pixelout<=1'b1;
37758: pixelout<=1'b1;
37759: pixelout<=1'b1;
37760: pixelout<=1'b1;
37761: pixelout<=1'b1;
37762: pixelout<=1'b1;
37763: pixelout<=1'b1;
37764: pixelout<=1'b1;
37765: pixelout<=1'b1;
37766: pixelout<=1'b1;
37767: pixelout<=1'b1;
37768: pixelout<=1'b1;
37769: pixelout<=1'b1;
37770: pixelout<=1'b1;
37771: pixelout<=1'b1;
37772: pixelout<=1'b1;
37773: pixelout<=1'b1;
37774: pixelout<=1'b1;
37775: pixelout<=1'b1;
37776: pixelout<=1'b1;
37777: pixelout<=1'b1;
37778: pixelout<=1'b1;
37779: pixelout<=1'b1;
37780: pixelout<=1'b1;
37781: pixelout<=1'b1;
37782: pixelout<=1'b1;
37783: pixelout<=1'b1;
37784: pixelout<=1'b1;
37785: pixelout<=1'b1;
37786: pixelout<=1'b1;
37787: pixelout<=1'b1;
37788: pixelout<=1'b1;
37789: pixelout<=1'b1;
37790: pixelout<=1'b1;
37791: pixelout<=1'b1;
37792: pixelout<=1'b1;
37793: pixelout<=1'b1;
37794: pixelout<=1'b1;
37795: pixelout<=1'b1;
37796: pixelout<=1'b1;
37797: pixelout<=1'b1;
37798: pixelout<=1'b1;
37799: pixelout<=1'b1;
37800: pixelout<=1'b1;
37801: pixelout<=1'b1;
37802: pixelout<=1'b1;
37803: pixelout<=1'b1;
37804: pixelout<=1'b1;
37805: pixelout<=1'b1;
37806: pixelout<=1'b1;
37807: pixelout<=1'b1;
37808: pixelout<=1'b1;
37809: pixelout<=1'b1;
37810: pixelout<=1'b1;
37811: pixelout<=1'b1;
37812: pixelout<=1'b1;
37813: pixelout<=1'b1;
37814: pixelout<=1'b1;
37815: pixelout<=1'b1;
37816: pixelout<=1'b1;
37817: pixelout<=1'b1;
37818: pixelout<=1'b1;
37819: pixelout<=1'b1;
37820: pixelout<=1'b1;
37821: pixelout<=1'b1;
37822: pixelout<=1'b1;
37823: pixelout<=1'b1;
37824: pixelout<=1'b1;
37825: pixelout<=1'b1;
37826: pixelout<=1'b1;
37827: pixelout<=1'b1;
37828: pixelout<=1'b1;
37829: pixelout<=1'b1;
37830: pixelout<=1'b1;
37831: pixelout<=1'b1;
37832: pixelout<=1'b1;
37833: pixelout<=1'b1;
37834: pixelout<=1'b1;
37835: pixelout<=1'b1;
37836: pixelout<=1'b1;
37837: pixelout<=1'b1;
37838: pixelout<=1'b1;
37839: pixelout<=1'b1;
37840: pixelout<=1'b1;
37841: pixelout<=1'b1;
37842: pixelout<=1'b1;
37843: pixelout<=1'b1;
37844: pixelout<=1'b1;
37845: pixelout<=1'b1;
37846: pixelout<=1'b1;
37847: pixelout<=1'b1;
37848: pixelout<=1'b1;
37849: pixelout<=1'b1;
37850: pixelout<=1'b1;
37851: pixelout<=1'b1;
37852: pixelout<=1'b1;
37853: pixelout<=1'b1;
37854: pixelout<=1'b1;
37855: pixelout<=1'b1;
37856: pixelout<=1'b1;
37857: pixelout<=1'b1;
37858: pixelout<=1'b1;
37859: pixelout<=1'b1;
37860: pixelout<=1'b1;
37861: pixelout<=1'b1;
37862: pixelout<=1'b1;
37863: pixelout<=1'b1;
37864: pixelout<=1'b1;
37865: pixelout<=1'b1;
37866: pixelout<=1'b1;
37867: pixelout<=1'b1;
37868: pixelout<=1'b1;
37869: pixelout<=1'b1;
37870: pixelout<=1'b1;
37871: pixelout<=1'b1;
37872: pixelout<=1'b1;
37873: pixelout<=1'b1;
37874: pixelout<=1'b1;
37875: pixelout<=1'b1;
37876: pixelout<=1'b1;
37877: pixelout<=1'b1;
37878: pixelout<=1'b1;
37879: pixelout<=1'b1;
37880: pixelout<=1'b1;
37881: pixelout<=1'b1;
37882: pixelout<=1'b1;
37883: pixelout<=1'b1;
37884: pixelout<=1'b1;
37885: pixelout<=1'b1;
37886: pixelout<=1'b1;
37887: pixelout<=1'b1;
37888: pixelout<=1'b1;
37889: pixelout<=1'b1;
37890: pixelout<=1'b1;
37891: pixelout<=1'b1;
37892: pixelout<=1'b1;
37893: pixelout<=1'b1;
37894: pixelout<=1'b1;
37895: pixelout<=1'b1;
37896: pixelout<=1'b1;
37897: pixelout<=1'b1;
37898: pixelout<=1'b1;
37899: pixelout<=1'b1;
37900: pixelout<=1'b1;
37901: pixelout<=1'b1;
37902: pixelout<=1'b1;
37903: pixelout<=1'b1;
37904: pixelout<=1'b1;
37905: pixelout<=1'b1;
37906: pixelout<=1'b1;
37907: pixelout<=1'b1;
37908: pixelout<=1'b1;
37909: pixelout<=1'b1;
37910: pixelout<=1'b1;
37911: pixelout<=1'b1;
37912: pixelout<=1'b1;
37913: pixelout<=1'b1;
37914: pixelout<=1'b1;
37915: pixelout<=1'b1;
37916: pixelout<=1'b1;
37917: pixelout<=1'b1;
37918: pixelout<=1'b1;
37919: pixelout<=1'b1;
37920: pixelout<=1'b1;
37921: pixelout<=1'b1;
37922: pixelout<=1'b1;
37923: pixelout<=1'b1;
37924: pixelout<=1'b1;
37925: pixelout<=1'b1;
37926: pixelout<=1'b1;
37927: pixelout<=1'b1;
37928: pixelout<=1'b1;
37929: pixelout<=1'b1;
37930: pixelout<=1'b1;
37931: pixelout<=1'b1;
37932: pixelout<=1'b1;
37933: pixelout<=1'b1;
37934: pixelout<=1'b1;
37935: pixelout<=1'b1;
37936: pixelout<=1'b1;
37937: pixelout<=1'b1;
37938: pixelout<=1'b1;
37939: pixelout<=1'b1;
37940: pixelout<=1'b1;
37941: pixelout<=1'b1;
37942: pixelout<=1'b1;
37943: pixelout<=1'b1;
37944: pixelout<=1'b1;
37945: pixelout<=1'b1;
37946: pixelout<=1'b1;
37947: pixelout<=1'b1;
37948: pixelout<=1'b1;
37949: pixelout<=1'b1;
37950: pixelout<=1'b1;
37951: pixelout<=1'b1;
37952: pixelout<=1'b1;
37953: pixelout<=1'b1;
37954: pixelout<=1'b1;
37955: pixelout<=1'b1;
37956: pixelout<=1'b1;
37957: pixelout<=1'b1;
37958: pixelout<=1'b1;
37959: pixelout<=1'b1;
37960: pixelout<=1'b1;
37961: pixelout<=1'b1;
37962: pixelout<=1'b1;
37963: pixelout<=1'b1;
37964: pixelout<=1'b1;
37965: pixelout<=1'b1;
37966: pixelout<=1'b1;
37967: pixelout<=1'b1;
37968: pixelout<=1'b1;
37969: pixelout<=1'b1;
37970: pixelout<=1'b1;
37971: pixelout<=1'b1;
37972: pixelout<=1'b1;
37973: pixelout<=1'b1;
37974: pixelout<=1'b1;
37975: pixelout<=1'b1;
37976: pixelout<=1'b1;
37977: pixelout<=1'b1;
37978: pixelout<=1'b1;
37979: pixelout<=1'b1;
37980: pixelout<=1'b1;
37981: pixelout<=1'b1;
37982: pixelout<=1'b1;
37983: pixelout<=1'b1;
37984: pixelout<=1'b1;
37985: pixelout<=1'b1;
37986: pixelout<=1'b1;
37987: pixelout<=1'b1;
37988: pixelout<=1'b1;
37989: pixelout<=1'b1;
37990: pixelout<=1'b1;
37991: pixelout<=1'b1;
37992: pixelout<=1'b1;
37993: pixelout<=1'b1;
37994: pixelout<=1'b1;
37995: pixelout<=1'b1;
37996: pixelout<=1'b1;
37997: pixelout<=1'b1;
37998: pixelout<=1'b1;
37999: pixelout<=1'b1;
38000: pixelout<=1'b1;
38001: pixelout<=1'b1;
38002: pixelout<=1'b1;
38003: pixelout<=1'b1;
38004: pixelout<=1'b1;
38005: pixelout<=1'b1;
38006: pixelout<=1'b1;
38007: pixelout<=1'b1;
38008: pixelout<=1'b1;
38009: pixelout<=1'b1;
38010: pixelout<=1'b1;
38011: pixelout<=1'b1;
38012: pixelout<=1'b1;
38013: pixelout<=1'b1;
38014: pixelout<=1'b1;
38015: pixelout<=1'b1;
38016: pixelout<=1'b1;
38017: pixelout<=1'b1;
38018: pixelout<=1'b1;
38019: pixelout<=1'b1;
38020: pixelout<=1'b1;
38021: pixelout<=1'b1;
38022: pixelout<=1'b1;
38023: pixelout<=1'b1;
38024: pixelout<=1'b1;
38025: pixelout<=1'b1;
38026: pixelout<=1'b1;
38027: pixelout<=1'b1;
38028: pixelout<=1'b1;
38029: pixelout<=1'b1;
38030: pixelout<=1'b1;
38031: pixelout<=1'b1;
38032: pixelout<=1'b1;
38033: pixelout<=1'b1;
38034: pixelout<=1'b1;
38035: pixelout<=1'b1;
38036: pixelout<=1'b1;
38037: pixelout<=1'b1;
38038: pixelout<=1'b1;
38039: pixelout<=1'b1;
38040: pixelout<=1'b1;
38041: pixelout<=1'b1;
38042: pixelout<=1'b1;
38043: pixelout<=1'b1;
38044: pixelout<=1'b1;
38045: pixelout<=1'b1;
38046: pixelout<=1'b1;
38047: pixelout<=1'b1;
38048: pixelout<=1'b1;
38049: pixelout<=1'b1;
38050: pixelout<=1'b1;
38051: pixelout<=1'b1;
38052: pixelout<=1'b1;
38053: pixelout<=1'b1;
38054: pixelout<=1'b1;
38055: pixelout<=1'b1;
38056: pixelout<=1'b1;
38057: pixelout<=1'b1;
38058: pixelout<=1'b1;
38059: pixelout<=1'b1;
38060: pixelout<=1'b1;
38061: pixelout<=1'b1;
38062: pixelout<=1'b1;
38063: pixelout<=1'b1;
38064: pixelout<=1'b1;
38065: pixelout<=1'b1;
38066: pixelout<=1'b1;
38067: pixelout<=1'b1;
38068: pixelout<=1'b1;
38069: pixelout<=1'b1;
38070: pixelout<=1'b1;
38071: pixelout<=1'b1;
38072: pixelout<=1'b1;
38073: pixelout<=1'b1;
38074: pixelout<=1'b1;
38075: pixelout<=1'b1;
38076: pixelout<=1'b1;
38077: pixelout<=1'b1;
38078: pixelout<=1'b1;
38079: pixelout<=1'b1;
38080: pixelout<=1'b1;
38081: pixelout<=1'b1;
38082: pixelout<=1'b1;
38083: pixelout<=1'b1;
38084: pixelout<=1'b1;
38085: pixelout<=1'b1;
38086: pixelout<=1'b1;
38087: pixelout<=1'b1;
38088: pixelout<=1'b1;
38089: pixelout<=1'b1;
38090: pixelout<=1'b1;
38091: pixelout<=1'b1;
38092: pixelout<=1'b1;
38093: pixelout<=1'b1;
38094: pixelout<=1'b1;
38095: pixelout<=1'b1;
38096: pixelout<=1'b1;
38097: pixelout<=1'b1;
38098: pixelout<=1'b1;
38099: pixelout<=1'b1;
38100: pixelout<=1'b1;
38101: pixelout<=1'b1;
38102: pixelout<=1'b1;
38103: pixelout<=1'b1;
38104: pixelout<=1'b1;
38105: pixelout<=1'b1;
38106: pixelout<=1'b1;
38107: pixelout<=1'b1;
38108: pixelout<=1'b1;
38109: pixelout<=1'b1;
38110: pixelout<=1'b1;
38111: pixelout<=1'b1;
38112: pixelout<=1'b1;
38113: pixelout<=1'b1;
38114: pixelout<=1'b1;
38115: pixelout<=1'b1;
38116: pixelout<=1'b1;
38117: pixelout<=1'b1;
38118: pixelout<=1'b1;
38119: pixelout<=1'b1;
38120: pixelout<=1'b1;
38121: pixelout<=1'b1;
38122: pixelout<=1'b1;
38123: pixelout<=1'b1;
38124: pixelout<=1'b1;
38125: pixelout<=1'b1;
38126: pixelout<=1'b1;
38127: pixelout<=1'b1;
38128: pixelout<=1'b1;
38129: pixelout<=1'b1;
38130: pixelout<=1'b1;
38131: pixelout<=1'b1;
38132: pixelout<=1'b1;
38133: pixelout<=1'b1;
38134: pixelout<=1'b1;
38135: pixelout<=1'b1;
38136: pixelout<=1'b1;
38137: pixelout<=1'b1;
38138: pixelout<=1'b1;
38139: pixelout<=1'b1;
38140: pixelout<=1'b1;
38141: pixelout<=1'b1;
38142: pixelout<=1'b1;
38143: pixelout<=1'b1;
38144: pixelout<=1'b1;
38145: pixelout<=1'b1;
38146: pixelout<=1'b1;
38147: pixelout<=1'b1;
38148: pixelout<=1'b1;
38149: pixelout<=1'b1;
38150: pixelout<=1'b1;
38151: pixelout<=1'b1;
38152: pixelout<=1'b1;
38153: pixelout<=1'b1;
38154: pixelout<=1'b1;
38155: pixelout<=1'b1;
38156: pixelout<=1'b1;
38157: pixelout<=1'b1;
38158: pixelout<=1'b1;
38159: pixelout<=1'b1;
38160: pixelout<=1'b1;
38161: pixelout<=1'b1;
38162: pixelout<=1'b1;
38163: pixelout<=1'b1;
38164: pixelout<=1'b1;
38165: pixelout<=1'b1;
38166: pixelout<=1'b1;
38167: pixelout<=1'b1;
38168: pixelout<=1'b1;
38169: pixelout<=1'b1;
38170: pixelout<=1'b1;
38171: pixelout<=1'b1;
38172: pixelout<=1'b1;
38173: pixelout<=1'b1;
38174: pixelout<=1'b1;
38175: pixelout<=1'b1;
38176: pixelout<=1'b1;
38177: pixelout<=1'b1;
38178: pixelout<=1'b1;
38179: pixelout<=1'b1;
38180: pixelout<=1'b1;
38181: pixelout<=1'b1;
38182: pixelout<=1'b1;
38183: pixelout<=1'b1;
38184: pixelout<=1'b1;
38185: pixelout<=1'b1;
38186: pixelout<=1'b1;
38187: pixelout<=1'b1;
38188: pixelout<=1'b1;
38189: pixelout<=1'b1;
38190: pixelout<=1'b1;
38191: pixelout<=1'b1;
38192: pixelout<=1'b1;
38193: pixelout<=1'b1;
38194: pixelout<=1'b1;
38195: pixelout<=1'b1;
38196: pixelout<=1'b1;
38197: pixelout<=1'b1;
38198: pixelout<=1'b1;
38199: pixelout<=1'b1;
38200: pixelout<=1'b1;
38201: pixelout<=1'b1;
38202: pixelout<=1'b1;
38203: pixelout<=1'b1;
38204: pixelout<=1'b1;
38205: pixelout<=1'b1;
38206: pixelout<=1'b1;
38207: pixelout<=1'b1;
38208: pixelout<=1'b1;
38209: pixelout<=1'b1;
38210: pixelout<=1'b1;
38211: pixelout<=1'b1;
38212: pixelout<=1'b1;
38213: pixelout<=1'b1;
38214: pixelout<=1'b1;
38215: pixelout<=1'b1;
38216: pixelout<=1'b1;
38217: pixelout<=1'b1;
38218: pixelout<=1'b1;
38219: pixelout<=1'b1;
38220: pixelout<=1'b1;
38221: pixelout<=1'b1;
38222: pixelout<=1'b1;
38223: pixelout<=1'b1;
38224: pixelout<=1'b1;
38225: pixelout<=1'b1;
38226: pixelout<=1'b1;
38227: pixelout<=1'b1;
38228: pixelout<=1'b1;
38229: pixelout<=1'b1;
38230: pixelout<=1'b1;
38231: pixelout<=1'b1;
38232: pixelout<=1'b1;
38233: pixelout<=1'b1;
38234: pixelout<=1'b1;
38235: pixelout<=1'b1;
38236: pixelout<=1'b1;
38237: pixelout<=1'b1;
38238: pixelout<=1'b1;
38239: pixelout<=1'b1;
38240: pixelout<=1'b1;
38241: pixelout<=1'b1;
38242: pixelout<=1'b1;
38243: pixelout<=1'b1;
38244: pixelout<=1'b1;
38245: pixelout<=1'b1;
38246: pixelout<=1'b1;
38247: pixelout<=1'b1;
38248: pixelout<=1'b1;
38249: pixelout<=1'b1;
38250: pixelout<=1'b1;
38251: pixelout<=1'b1;
38252: pixelout<=1'b1;
38253: pixelout<=1'b1;
38254: pixelout<=1'b1;
38255: pixelout<=1'b1;
38256: pixelout<=1'b1;
38257: pixelout<=1'b1;
38258: pixelout<=1'b1;
38259: pixelout<=1'b1;
38260: pixelout<=1'b1;
38261: pixelout<=1'b1;
38262: pixelout<=1'b1;
38263: pixelout<=1'b1;
38264: pixelout<=1'b1;
38265: pixelout<=1'b1;
38266: pixelout<=1'b1;
38267: pixelout<=1'b1;
38268: pixelout<=1'b1;
38269: pixelout<=1'b1;
38270: pixelout<=1'b1;
38271: pixelout<=1'b1;
38272: pixelout<=1'b1;
38273: pixelout<=1'b1;
38274: pixelout<=1'b1;
38275: pixelout<=1'b1;
38276: pixelout<=1'b1;
38277: pixelout<=1'b1;
38278: pixelout<=1'b1;
38279: pixelout<=1'b1;
38280: pixelout<=1'b1;
38281: pixelout<=1'b1;
38282: pixelout<=1'b1;
38283: pixelout<=1'b1;
38284: pixelout<=1'b1;
38285: pixelout<=1'b1;
38286: pixelout<=1'b1;
38287: pixelout<=1'b1;
38288: pixelout<=1'b1;
38289: pixelout<=1'b1;
38290: pixelout<=1'b1;
38291: pixelout<=1'b1;
38292: pixelout<=1'b1;
38293: pixelout<=1'b1;
38294: pixelout<=1'b1;
38295: pixelout<=1'b1;
38296: pixelout<=1'b1;
38297: pixelout<=1'b1;
38298: pixelout<=1'b1;
38299: pixelout<=1'b1;
38300: pixelout<=1'b1;
38301: pixelout<=1'b1;
38302: pixelout<=1'b1;
38303: pixelout<=1'b1;
38304: pixelout<=1'b1;
38305: pixelout<=1'b1;
38306: pixelout<=1'b1;
38307: pixelout<=1'b1;
38308: pixelout<=1'b1;
38309: pixelout<=1'b1;
38310: pixelout<=1'b1;
38311: pixelout<=1'b1;
38312: pixelout<=1'b1;
38313: pixelout<=1'b1;
38314: pixelout<=1'b1;
38315: pixelout<=1'b1;
38316: pixelout<=1'b1;
38317: pixelout<=1'b1;
38318: pixelout<=1'b1;
38319: pixelout<=1'b1;
38320: pixelout<=1'b1;
38321: pixelout<=1'b1;
38322: pixelout<=1'b1;
38323: pixelout<=1'b1;
38324: pixelout<=1'b1;
38325: pixelout<=1'b1;
38326: pixelout<=1'b1;
38327: pixelout<=1'b1;
38328: pixelout<=1'b1;
38329: pixelout<=1'b1;
38330: pixelout<=1'b1;
38331: pixelout<=1'b1;
38332: pixelout<=1'b1;
38333: pixelout<=1'b1;
38334: pixelout<=1'b1;
38335: pixelout<=1'b1;
38336: pixelout<=1'b1;
38337: pixelout<=1'b1;
38338: pixelout<=1'b1;
38339: pixelout<=1'b1;
38340: pixelout<=1'b1;
38341: pixelout<=1'b1;
38342: pixelout<=1'b1;
38343: pixelout<=1'b1;
38344: pixelout<=1'b1;
38345: pixelout<=1'b1;
38346: pixelout<=1'b1;
38347: pixelout<=1'b1;
38348: pixelout<=1'b1;
38349: pixelout<=1'b1;
38350: pixelout<=1'b1;
38351: pixelout<=1'b1;
38352: pixelout<=1'b1;
38353: pixelout<=1'b1;
38354: pixelout<=1'b1;
38355: pixelout<=1'b1;
38356: pixelout<=1'b1;
38357: pixelout<=1'b1;
38358: pixelout<=1'b1;
38359: pixelout<=1'b1;
38360: pixelout<=1'b1;
38361: pixelout<=1'b1;
38362: pixelout<=1'b1;
38363: pixelout<=1'b1;
38364: pixelout<=1'b1;
38365: pixelout<=1'b1;
38366: pixelout<=1'b1;
38367: pixelout<=1'b1;
38368: pixelout<=1'b1;
38369: pixelout<=1'b1;
38370: pixelout<=1'b1;
38371: pixelout<=1'b1;
38372: pixelout<=1'b1;
38373: pixelout<=1'b1;
38374: pixelout<=1'b1;
38375: pixelout<=1'b1;
38376: pixelout<=1'b1;
38377: pixelout<=1'b1;
38378: pixelout<=1'b1;
38379: pixelout<=1'b1;
38380: pixelout<=1'b1;
38381: pixelout<=1'b1;
38382: pixelout<=1'b1;
38383: pixelout<=1'b1;
38384: pixelout<=1'b1;
38385: pixelout<=1'b1;
38386: pixelout<=1'b1;
38387: pixelout<=1'b1;
38388: pixelout<=1'b1;
38389: pixelout<=1'b1;
38390: pixelout<=1'b1;
38391: pixelout<=1'b1;
38392: pixelout<=1'b1;
38393: pixelout<=1'b1;
38394: pixelout<=1'b1;
38395: pixelout<=1'b1;
38396: pixelout<=1'b1;
38397: pixelout<=1'b1;
38398: pixelout<=1'b1;
38399: pixelout<=1'b1;
default : ; 
endcase
end
endmodule