module fakeramlol (input clk, input[15:0] n, output pixelout)

always_ff @ (posedge clk)
begin
case (n)
	0 : 1;
	1 : 1;
	2 : 1;
	3 : 1;
	4 : 1;
	5 : 1;
	6 : 1;
	7 : 1;
	8 : 1;
	9 : 1;
	10 : 1;
	11 : 1;
	12 : 1;
	13 : 1;
	14 : 1;
	15 : 1;
	16 : 1;
	17 : 1;
	18 : 1;
	19 : 1;
	20 : 1;
	21 : 1;
	22 : 1;
	23 : 1;
	24 : 1;
	25 : 1;
	26 : 1;
	27 : 1;
	28 : 1;
	29 : 1;
	30 : 1;
	31 : 1;
	32 : 1;
	33 : 1;
	34 : 1;
	35 : 1;
	36 : 1;
	37 : 1;
	38 : 1;
	39 : 1;
	40 : 1;
	41 : 1;
	42 : 1;
	43 : 1;
	44 : 1;
	45 : 1;
	46 : 1;
	47 : 1;
	48 : 1;
	49 : 1;
	50 : 1;
	51 : 1;
	52 : 1;
	53 : 1;
	54 : 1;
	55 : 1;
	56 : 1;
	57 : 1;
	58 : 1;
	59 : 1;
	60 : 1;
	61 : 1;
	62 : 1;
	63 : 1;
	64 : 1;
	65 : 1;
	66 : 1;
	67 : 1;
	68 : 1;
	69 : 1;
	70 : 1;
	71 : 1;
	72 : 1;
	73 : 1;
	74 : 1;
	75 : 1;
	76 : 1;
	77 : 1;
	78 : 1;
	79 : 1;
	80 : 1;
	81 : 1;
	82 : 1;
	83 : 1;
	84 : 1;
	85 : 1;
	86 : 1;
	87 : 1;
	88 : 1;
	89 : 1;
	90 : 1;
	91 : 1;
	92 : 1;
	93 : 1;
	94 : 1;
	95 : 1;
	96 : 1;
	97 : 1;
	98 : 1;
	99 : 1;
	100 : 1;
	101 : 1;
	102 : 1;
	103 : 1;
	104 : 1;
	105 : 1;
	106 : 1;
	107 : 1;
	108 : 1;
	109 : 1;
	110 : 1;
	111 : 1;
	112 : 1;
	113 : 1;
	114 : 1;
	115 : 1;
	116 : 1;
	117 : 1;
	118 : 1;
	119 : 1;
	120 : 1;
	121 : 1;
	122 : 1;
	123 : 1;
	124 : 1;
	125 : 1;
	126 : 1;
	127 : 1;
	128 : 1;
	129 : 1;
	130 : 1;
	131 : 1;
	132 : 1;
	133 : 1;
	134 : 1;
	135 : 1;
	136 : 1;
	137 : 1;
	138 : 1;
	139 : 1;
	140 : 1;
	141 : 1;
	142 : 1;
	143 : 1;
	144 : 1;
	145 : 1;
	146 : 1;
	147 : 1;
	148 : 1;
	149 : 1;
	150 : 1;
	151 : 1;
	152 : 1;
	153 : 1;
	154 : 1;
	155 : 1;
	156 : 1;
	157 : 1;
	158 : 1;
	159 : 1;
	160 : 1;
	161 : 1;
	162 : 1;
	163 : 1;
	164 : 1;
	165 : 1;
	166 : 1;
	167 : 1;
	168 : 1;
	169 : 1;
	170 : 1;
	171 : 1;
	172 : 1;
	173 : 1;
	174 : 1;
	175 : 1;
	176 : 1;
	177 : 1;
	178 : 1;
	179 : 1;
	180 : 1;
	181 : 1;
	182 : 1;
	183 : 1;
	184 : 1;
	185 : 1;
	186 : 1;
	187 : 1;
	188 : 1;
	189 : 1;
	190 : 1;
	191 : 1;
	192 : 1;
	193 : 1;
	194 : 1;
	195 : 1;
	196 : 1;
	197 : 1;
	198 : 1;
	199 : 1;
	200 : 1;
	201 : 1;
	202 : 1;
	203 : 1;
	204 : 1;
	205 : 1;
	206 : 1;
	207 : 1;
	208 : 1;
	209 : 1;
	210 : 1;
	211 : 1;
	212 : 1;
	213 : 1;
	214 : 1;
	215 : 1;
	216 : 1;
	217 : 1;
	218 : 1;
	219 : 1;
	220 : 1;
	221 : 1;
	222 : 1;
	223 : 1;
	224 : 1;
	225 : 1;
	226 : 1;
	227 : 1;
	228 : 1;
	229 : 1;
	230 : 1;
	231 : 1;
	232 : 1;
	233 : 1;
	234 : 1;
	235 : 1;
	236 : 1;
	237 : 1;
	238 : 1;
	239 : 1;
	240 : 1;
	241 : 1;
	242 : 1;
	243 : 1;
	244 : 1;
	245 : 1;
	246 : 1;
	247 : 1;
	248 : 1;
	249 : 1;
	250 : 1;
	251 : 1;
	252 : 1;
	253 : 1;
	254 : 1;
	255 : 1;
	256 : 1;
	257 : 1;
	258 : 1;
	259 : 1;
	260 : 1;
	261 : 1;
	262 : 1;
	263 : 1;
	264 : 1;
	265 : 1;
	266 : 1;
	267 : 1;
	268 : 1;
	269 : 1;
	270 : 1;
	271 : 1;
	272 : 1;
	273 : 1;
	274 : 1;
	275 : 1;
	276 : 1;
	277 : 1;
	278 : 1;
	279 : 1;
	280 : 1;
	281 : 1;
	282 : 1;
	283 : 1;
	284 : 1;
	285 : 1;
	286 : 1;
	287 : 1;
	288 : 1;
	289 : 1;
	290 : 1;
	291 : 1;
	292 : 1;
	293 : 1;
	294 : 1;
	295 : 1;
	296 : 1;
	297 : 1;
	298 : 1;
	299 : 1;
	300 : 1;
	301 : 1;
	302 : 1;
	303 : 1;
	304 : 1;
	305 : 1;
	306 : 1;
	307 : 1;
	308 : 1;
	309 : 1;
	310 : 1;
	311 : 1;
	312 : 1;
	313 : 1;
	314 : 1;
	315 : 1;
	316 : 1;
	317 : 1;
	318 : 1;
	319 : 1;
	320 : 1;
	321 : 1;
	322 : 1;
	323 : 1;
	324 : 1;
	325 : 1;
	326 : 1;
	327 : 1;
	328 : 1;
	329 : 1;
	330 : 1;
	331 : 1;
	332 : 1;
	333 : 1;
	334 : 1;
	335 : 1;
	336 : 1;
	337 : 1;
	338 : 1;
	339 : 1;
	340 : 1;
	341 : 1;
	342 : 1;
	343 : 1;
	344 : 1;
	345 : 1;
	346 : 1;
	347 : 1;
	348 : 1;
	349 : 1;
	350 : 1;
	351 : 1;
	352 : 1;
	353 : 1;
	354 : 1;
	355 : 1;
	356 : 1;
	357 : 1;
	358 : 1;
	359 : 1;
	360 : 1;
	361 : 1;
	362 : 1;
	363 : 1;
	364 : 1;
	365 : 1;
	366 : 1;
	367 : 1;
	368 : 1;
	369 : 1;
	370 : 1;
	371 : 1;
	372 : 1;
	373 : 1;
	374 : 1;
	375 : 1;
	376 : 1;
	377 : 1;
	378 : 1;
	379 : 1;
	380 : 1;
	381 : 1;
	382 : 1;
	383 : 1;
	384 : 1;
	385 : 1;
	386 : 1;
	387 : 1;
	388 : 1;
	389 : 1;
	390 : 1;
	391 : 1;
	392 : 1;
	393 : 1;
	394 : 1;
	395 : 1;
	396 : 1;
	397 : 1;
	398 : 1;
	399 : 1;
	400 : 1;
	401 : 1;
	402 : 1;
	403 : 1;
	404 : 1;
	405 : 1;
	406 : 1;
	407 : 1;
	408 : 1;
	409 : 1;
	410 : 1;
	411 : 1;
	412 : 1;
	413 : 1;
	414 : 1;
	415 : 1;
	416 : 1;
	417 : 1;
	418 : 1;
	419 : 1;
	420 : 1;
	421 : 1;
	422 : 1;
	423 : 1;
	424 : 1;
	425 : 1;
	426 : 1;
	427 : 1;
	428 : 1;
	429 : 1;
	430 : 1;
	431 : 1;
	432 : 1;
	433 : 1;
	434 : 1;
	435 : 1;
	436 : 1;
	437 : 1;
	438 : 1;
	439 : 1;
	440 : 1;
	441 : 1;
	442 : 1;
	443 : 1;
	444 : 1;
	445 : 1;
	446 : 1;
	447 : 1;
	448 : 1;
	449 : 1;
	450 : 1;
	451 : 1;
	452 : 1;
	453 : 1;
	454 : 1;
	455 : 1;
	456 : 1;
	457 : 1;
	458 : 1;
	459 : 1;
	460 : 1;
	461 : 1;
	462 : 1;
	463 : 1;
	464 : 1;
	465 : 1;
	466 : 1;
	467 : 1;
	468 : 1;
	469 : 1;
	470 : 1;
	471 : 1;
	472 : 1;
	473 : 1;
	474 : 1;
	475 : 1;
	476 : 1;
	477 : 1;
	478 : 1;
	479 : 1;
	480 : 1;
	481 : 1;
	482 : 1;
	483 : 1;
	484 : 1;
	485 : 1;
	486 : 1;
	487 : 1;
	488 : 1;
	489 : 1;
	490 : 1;
	491 : 1;
	492 : 1;
	493 : 1;
	494 : 1;
	495 : 1;
	496 : 1;
	497 : 1;
	498 : 1;
	499 : 1;
	500 : 1;
	501 : 1;
	502 : 1;
	503 : 1;
	504 : 1;
	505 : 1;
	506 : 1;
	507 : 1;
	508 : 1;
	509 : 1;
	510 : 1;
	511 : 1;
	512 : 1;
	513 : 1;
	514 : 1;
	515 : 1;
	516 : 1;
	517 : 1;
	518 : 1;
	519 : 1;
	520 : 1;
	521 : 1;
	522 : 1;
	523 : 1;
	524 : 1;
	525 : 1;
	526 : 1;
	527 : 1;
	528 : 1;
	529 : 1;
	530 : 1;
	531 : 1;
	532 : 1;
	533 : 1;
	534 : 1;
	535 : 1;
	536 : 1;
	537 : 1;
	538 : 1;
	539 : 1;
	540 : 1;
	541 : 1;
	542 : 1;
	543 : 1;
	544 : 1;
	545 : 1;
	546 : 1;
	547 : 1;
	548 : 1;
	549 : 1;
	550 : 1;
	551 : 1;
	552 : 1;
	553 : 1;
	554 : 1;
	555 : 1;
	556 : 1;
	557 : 1;
	558 : 1;
	559 : 1;
	560 : 1;
	561 : 1;
	562 : 1;
	563 : 1;
	564 : 1;
	565 : 1;
	566 : 1;
	567 : 1;
	568 : 1;
	569 : 1;
	570 : 1;
	571 : 1;
	572 : 1;
	573 : 1;
	574 : 1;
	575 : 1;
	576 : 1;
	577 : 1;
	578 : 1;
	579 : 1;
	580 : 1;
	581 : 1;
	582 : 1;
	583 : 1;
	584 : 1;
	585 : 1;
	586 : 1;
	587 : 1;
	588 : 1;
	589 : 1;
	590 : 1;
	591 : 1;
	592 : 1;
	593 : 1;
	594 : 1;
	595 : 1;
	596 : 1;
	597 : 1;
	598 : 1;
	599 : 1;
	600 : 1;
	601 : 1;
	602 : 1;
	603 : 1;
	604 : 1;
	605 : 1;
	606 : 1;
	607 : 1;
	608 : 1;
	609 : 1;
	610 : 1;
	611 : 1;
	612 : 1;
	613 : 1;
	614 : 1;
	615 : 1;
	616 : 1;
	617 : 1;
	618 : 1;
	619 : 1;
	620 : 1;
	621 : 1;
	622 : 1;
	623 : 1;
	624 : 1;
	625 : 1;
	626 : 1;
	627 : 1;
	628 : 1;
	629 : 1;
	630 : 1;
	631 : 1;
	632 : 1;
	633 : 1;
	634 : 1;
	635 : 1;
	636 : 1;
	637 : 1;
	638 : 1;
	639 : 1;
	640 : 1;
	641 : 1;
	642 : 1;
	643 : 1;
	644 : 1;
	645 : 1;
	646 : 1;
	647 : 1;
	648 : 1;
	649 : 1;
	650 : 1;
	651 : 1;
	652 : 1;
	653 : 1;
	654 : 1;
	655 : 1;
	656 : 1;
	657 : 1;
	658 : 1;
	659 : 1;
	660 : 1;
	661 : 1;
	662 : 1;
	663 : 1;
	664 : 1;
	665 : 1;
	666 : 1;
	667 : 1;
	668 : 1;
	669 : 1;
	670 : 1;
	671 : 1;
	672 : 1;
	673 : 1;
	674 : 1;
	675 : 1;
	676 : 1;
	677 : 1;
	678 : 1;
	679 : 1;
	680 : 1;
	681 : 1;
	682 : 1;
	683 : 1;
	684 : 1;
	685 : 1;
	686 : 1;
	687 : 1;
	688 : 1;
	689 : 1;
	690 : 1;
	691 : 1;
	692 : 1;
	693 : 1;
	694 : 1;
	695 : 1;
	696 : 1;
	697 : 1;
	698 : 1;
	699 : 1;
	700 : 1;
	701 : 1;
	702 : 1;
	703 : 1;
	704 : 1;
	705 : 1;
	706 : 1;
	707 : 1;
	708 : 1;
	709 : 1;
	710 : 1;
	711 : 1;
	712 : 1;
	713 : 1;
	714 : 1;
	715 : 1;
	716 : 1;
	717 : 1;
	718 : 1;
	719 : 1;
	720 : 1;
	721 : 1;
	722 : 1;
	723 : 1;
	724 : 1;
	725 : 1;
	726 : 1;
	727 : 1;
	728 : 1;
	729 : 1;
	730 : 1;
	731 : 1;
	732 : 1;
	733 : 1;
	734 : 1;
	735 : 1;
	736 : 1;
	737 : 1;
	738 : 1;
	739 : 1;
	740 : 1;
	741 : 1;
	742 : 1;
	743 : 1;
	744 : 1;
	745 : 1;
	746 : 1;
	747 : 1;
	748 : 1;
	749 : 1;
	750 : 1;
	751 : 1;
	752 : 1;
	753 : 1;
	754 : 1;
	755 : 1;
	756 : 1;
	757 : 1;
	758 : 1;
	759 : 1;
	760 : 1;
	761 : 1;
	762 : 1;
	763 : 1;
	764 : 1;
	765 : 1;
	766 : 1;
	767 : 1;
	768 : 1;
	769 : 1;
	770 : 1;
	771 : 1;
	772 : 1;
	773 : 1;
	774 : 1;
	775 : 1;
	776 : 1;
	777 : 1;
	778 : 1;
	779 : 1;
	780 : 1;
	781 : 1;
	782 : 1;
	783 : 1;
	784 : 1;
	785 : 1;
	786 : 1;
	787 : 1;
	788 : 1;
	789 : 1;
	790 : 1;
	791 : 1;
	792 : 1;
	793 : 1;
	794 : 1;
	795 : 1;
	796 : 1;
	797 : 1;
	798 : 1;
	799 : 1;
	800 : 1;
	801 : 1;
	802 : 1;
	803 : 1;
	804 : 1;
	805 : 1;
	806 : 1;
	807 : 1;
	808 : 1;
	809 : 1;
	810 : 1;
	811 : 1;
	812 : 1;
	813 : 1;
	814 : 1;
	815 : 1;
	816 : 1;
	817 : 1;
	818 : 1;
	819 : 1;
	820 : 1;
	821 : 1;
	822 : 1;
	823 : 1;
	824 : 1;
	825 : 1;
	826 : 1;
	827 : 1;
	828 : 1;
	829 : 1;
	830 : 1;
	831 : 1;
	832 : 1;
	833 : 1;
	834 : 1;
	835 : 1;
	836 : 1;
	837 : 1;
	838 : 1;
	839 : 1;
	840 : 1;
	841 : 1;
	842 : 1;
	843 : 1;
	844 : 1;
	845 : 1;
	846 : 1;
	847 : 1;
	848 : 1;
	849 : 1;
	850 : 1;
	851 : 1;
	852 : 1;
	853 : 1;
	854 : 1;
	855 : 1;
	856 : 1;
	857 : 1;
	858 : 1;
	859 : 1;
	860 : 1;
	861 : 1;
	862 : 1;
	863 : 1;
	864 : 1;
	865 : 1;
	866 : 1;
	867 : 1;
	868 : 1;
	869 : 1;
	870 : 1;
	871 : 1;
	872 : 1;
	873 : 1;
	874 : 1;
	875 : 1;
	876 : 1;
	877 : 1;
	878 : 1;
	879 : 1;
	880 : 1;
	881 : 1;
	882 : 1;
	883 : 1;
	884 : 1;
	885 : 1;
	886 : 1;
	887 : 1;
	888 : 1;
	889 : 1;
	890 : 1;
	891 : 1;
	892 : 1;
	893 : 1;
	894 : 1;
	895 : 1;
	896 : 1;
	897 : 1;
	898 : 1;
	899 : 1;
	900 : 1;
	901 : 1;
	902 : 1;
	903 : 1;
	904 : 1;
	905 : 1;
	906 : 1;
	907 : 1;
	908 : 1;
	909 : 1;
	910 : 1;
	911 : 1;
	912 : 1;
	913 : 1;
	914 : 1;
	915 : 1;
	916 : 1;
	917 : 1;
	918 : 1;
	919 : 1;
	920 : 1;
	921 : 1;
	922 : 1;
	923 : 1;
	924 : 1;
	925 : 1;
	926 : 1;
	927 : 1;
	928 : 1;
	929 : 1;
	930 : 1;
	931 : 1;
	932 : 1;
	933 : 1;
	934 : 1;
	935 : 1;
	936 : 1;
	937 : 1;
	938 : 1;
	939 : 1;
	940 : 1;
	941 : 1;
	942 : 1;
	943 : 1;
	944 : 1;
	945 : 1;
	946 : 1;
	947 : 1;
	948 : 1;
	949 : 1;
	950 : 1;
	951 : 1;
	952 : 1;
	953 : 1;
	954 : 1;
	955 : 1;
	956 : 1;
	957 : 1;
	958 : 1;
	959 : 1;
	960 : 1;
	961 : 1;
	962 : 1;
	963 : 1;
	964 : 1;
	965 : 1;
	966 : 1;
	967 : 1;
	968 : 1;
	969 : 1;
	970 : 1;
	971 : 1;
	972 : 1;
	973 : 1;
	974 : 1;
	975 : 1;
	976 : 1;
	977 : 1;
	978 : 1;
	979 : 1;
	980 : 1;
	981 : 1;
	982 : 1;
	983 : 1;
	984 : 1;
	985 : 1;
	986 : 1;
	987 : 1;
	988 : 1;
	989 : 1;
	990 : 1;
	991 : 1;
	992 : 1;
	993 : 1;
	994 : 1;
	995 : 1;
	996 : 1;
	997 : 1;
	998 : 1;
	999 : 1;
	1000 : 1;
	1001 : 1;
	1002 : 1;
	1003 : 1;
	1004 : 1;
	1005 : 1;
	1006 : 1;
	1007 : 1;
	1008 : 1;
	1009 : 1;
	1010 : 1;
	1011 : 1;
	1012 : 1;
	1013 : 1;
	1014 : 1;
	1015 : 1;
	1016 : 1;
	1017 : 1;
	1018 : 1;
	1019 : 1;
	1020 : 1;
	1021 : 1;
	1022 : 1;
	1023 : 1;
	1024 : 1;
	1025 : 1;
	1026 : 1;
	1027 : 1;
	1028 : 1;
	1029 : 1;
	1030 : 1;
	1031 : 1;
	1032 : 1;
	1033 : 1;
	1034 : 1;
	1035 : 1;
	1036 : 1;
	1037 : 1;
	1038 : 1;
	1039 : 1;
	1040 : 1;
	1041 : 1;
	1042 : 1;
	1043 : 1;
	1044 : 1;
	1045 : 1;
	1046 : 1;
	1047 : 1;
	1048 : 1;
	1049 : 1;
	1050 : 1;
	1051 : 1;
	1052 : 1;
	1053 : 1;
	1054 : 1;
	1055 : 1;
	1056 : 1;
	1057 : 1;
	1058 : 1;
	1059 : 1;
	1060 : 1;
	1061 : 1;
	1062 : 1;
	1063 : 1;
	1064 : 1;
	1065 : 1;
	1066 : 1;
	1067 : 1;
	1068 : 1;
	1069 : 1;
	1070 : 1;
	1071 : 1;
	1072 : 1;
	1073 : 1;
	1074 : 1;
	1075 : 1;
	1076 : 1;
	1077 : 1;
	1078 : 1;
	1079 : 1;
	1080 : 1;
	1081 : 1;
	1082 : 1;
	1083 : 1;
	1084 : 1;
	1085 : 1;
	1086 : 1;
	1087 : 1;
	1088 : 1;
	1089 : 1;
	1090 : 1;
	1091 : 1;
	1092 : 1;
	1093 : 1;
	1094 : 1;
	1095 : 1;
	1096 : 1;
	1097 : 1;
	1098 : 1;
	1099 : 1;
	1100 : 1;
	1101 : 1;
	1102 : 1;
	1103 : 1;
	1104 : 1;
	1105 : 1;
	1106 : 1;
	1107 : 1;
	1108 : 1;
	1109 : 1;
	1110 : 1;
	1111 : 1;
	1112 : 1;
	1113 : 1;
	1114 : 1;
	1115 : 1;
	1116 : 1;
	1117 : 1;
	1118 : 1;
	1119 : 1;
	1120 : 1;
	1121 : 1;
	1122 : 1;
	1123 : 1;
	1124 : 1;
	1125 : 1;
	1126 : 1;
	1127 : 1;
	1128 : 1;
	1129 : 1;
	1130 : 1;
	1131 : 1;
	1132 : 1;
	1133 : 1;
	1134 : 1;
	1135 : 1;
	1136 : 1;
	1137 : 1;
	1138 : 1;
	1139 : 1;
	1140 : 1;
	1141 : 1;
	1142 : 1;
	1143 : 1;
	1144 : 1;
	1145 : 1;
	1146 : 1;
	1147 : 1;
	1148 : 1;
	1149 : 1;
	1150 : 1;
	1151 : 1;
	1152 : 1;
	1153 : 1;
	1154 : 1;
	1155 : 1;
	1156 : 1;
	1157 : 1;
	1158 : 1;
	1159 : 1;
	1160 : 1;
	1161 : 1;
	1162 : 1;
	1163 : 1;
	1164 : 1;
	1165 : 1;
	1166 : 1;
	1167 : 1;
	1168 : 1;
	1169 : 1;
	1170 : 1;
	1171 : 1;
	1172 : 1;
	1173 : 1;
	1174 : 1;
	1175 : 1;
	1176 : 1;
	1177 : 1;
	1178 : 1;
	1179 : 1;
	1180 : 1;
	1181 : 1;
	1182 : 1;
	1183 : 1;
	1184 : 1;
	1185 : 1;
	1186 : 1;
	1187 : 1;
	1188 : 1;
	1189 : 1;
	1190 : 1;
	1191 : 1;
	1192 : 1;
	1193 : 1;
	1194 : 1;
	1195 : 1;
	1196 : 1;
	1197 : 1;
	1198 : 1;
	1199 : 1;
	1200 : 1;
	1201 : 1;
	1202 : 1;
	1203 : 1;
	1204 : 1;
	1205 : 1;
	1206 : 1;
	1207 : 1;
	1208 : 1;
	1209 : 1;
	1210 : 1;
	1211 : 1;
	1212 : 1;
	1213 : 1;
	1214 : 1;
	1215 : 1;
	1216 : 1;
	1217 : 1;
	1218 : 1;
	1219 : 1;
	1220 : 1;
	1221 : 1;
	1222 : 1;
	1223 : 1;
	1224 : 1;
	1225 : 1;
	1226 : 1;
	1227 : 1;
	1228 : 1;
	1229 : 1;
	1230 : 1;
	1231 : 1;
	1232 : 1;
	1233 : 1;
	1234 : 1;
	1235 : 1;
	1236 : 1;
	1237 : 1;
	1238 : 1;
	1239 : 1;
	1240 : 1;
	1241 : 1;
	1242 : 1;
	1243 : 1;
	1244 : 1;
	1245 : 1;
	1246 : 1;
	1247 : 1;
	1248 : 1;
	1249 : 1;
	1250 : 1;
	1251 : 1;
	1252 : 1;
	1253 : 1;
	1254 : 1;
	1255 : 1;
	1256 : 1;
	1257 : 1;
	1258 : 1;
	1259 : 1;
	1260 : 1;
	1261 : 1;
	1262 : 1;
	1263 : 1;
	1264 : 1;
	1265 : 1;
	1266 : 1;
	1267 : 1;
	1268 : 1;
	1269 : 1;
	1270 : 1;
	1271 : 1;
	1272 : 1;
	1273 : 1;
	1274 : 1;
	1275 : 1;
	1276 : 1;
	1277 : 1;
	1278 : 1;
	1279 : 1;
	1280 : 1;
	1281 : 1;
	1282 : 1;
	1283 : 1;
	1284 : 1;
	1285 : 1;
	1286 : 1;
	1287 : 1;
	1288 : 1;
	1289 : 1;
	1290 : 1;
	1291 : 1;
	1292 : 1;
	1293 : 1;
	1294 : 1;
	1295 : 1;
	1296 : 1;
	1297 : 1;
	1298 : 1;
	1299 : 1;
	1300 : 1;
	1301 : 1;
	1302 : 1;
	1303 : 1;
	1304 : 1;
	1305 : 1;
	1306 : 1;
	1307 : 1;
	1308 : 1;
	1309 : 1;
	1310 : 1;
	1311 : 1;
	1312 : 1;
	1313 : 1;
	1314 : 1;
	1315 : 1;
	1316 : 1;
	1317 : 1;
	1318 : 1;
	1319 : 1;
	1320 : 1;
	1321 : 1;
	1322 : 1;
	1323 : 1;
	1324 : 1;
	1325 : 1;
	1326 : 1;
	1327 : 1;
	1328 : 1;
	1329 : 1;
	1330 : 1;
	1331 : 1;
	1332 : 1;
	1333 : 1;
	1334 : 1;
	1335 : 1;
	1336 : 1;
	1337 : 1;
	1338 : 1;
	1339 : 1;
	1340 : 1;
	1341 : 1;
	1342 : 1;
	1343 : 1;
	1344 : 1;
	1345 : 1;
	1346 : 1;
	1347 : 1;
	1348 : 1;
	1349 : 1;
	1350 : 1;
	1351 : 1;
	1352 : 1;
	1353 : 1;
	1354 : 1;
	1355 : 1;
	1356 : 1;
	1357 : 1;
	1358 : 1;
	1359 : 1;
	1360 : 1;
	1361 : 1;
	1362 : 1;
	1363 : 1;
	1364 : 1;
	1365 : 1;
	1366 : 1;
	1367 : 1;
	1368 : 1;
	1369 : 1;
	1370 : 1;
	1371 : 1;
	1372 : 1;
	1373 : 1;
	1374 : 1;
	1375 : 1;
	1376 : 1;
	1377 : 1;
	1378 : 1;
	1379 : 1;
	1380 : 1;
	1381 : 1;
	1382 : 1;
	1383 : 1;
	1384 : 1;
	1385 : 1;
	1386 : 1;
	1387 : 1;
	1388 : 1;
	1389 : 1;
	1390 : 1;
	1391 : 1;
	1392 : 1;
	1393 : 1;
	1394 : 1;
	1395 : 1;
	1396 : 1;
	1397 : 1;
	1398 : 1;
	1399 : 1;
	1400 : 1;
	1401 : 1;
	1402 : 1;
	1403 : 1;
	1404 : 1;
	1405 : 1;
	1406 : 1;
	1407 : 1;
	1408 : 1;
	1409 : 1;
	1410 : 1;
	1411 : 1;
	1412 : 1;
	1413 : 1;
	1414 : 1;
	1415 : 1;
	1416 : 1;
	1417 : 1;
	1418 : 1;
	1419 : 1;
	1420 : 1;
	1421 : 1;
	1422 : 1;
	1423 : 1;
	1424 : 1;
	1425 : 1;
	1426 : 1;
	1427 : 1;
	1428 : 1;
	1429 : 1;
	1430 : 1;
	1431 : 1;
	1432 : 1;
	1433 : 1;
	1434 : 1;
	1435 : 1;
	1436 : 1;
	1437 : 1;
	1438 : 1;
	1439 : 1;
	1440 : 1;
	1441 : 1;
	1442 : 1;
	1443 : 1;
	1444 : 1;
	1445 : 1;
	1446 : 1;
	1447 : 1;
	1448 : 1;
	1449 : 1;
	1450 : 1;
	1451 : 1;
	1452 : 1;
	1453 : 1;
	1454 : 1;
	1455 : 1;
	1456 : 1;
	1457 : 1;
	1458 : 1;
	1459 : 1;
	1460 : 1;
	1461 : 1;
	1462 : 1;
	1463 : 1;
	1464 : 1;
	1465 : 1;
	1466 : 1;
	1467 : 1;
	1468 : 1;
	1469 : 1;
	1470 : 1;
	1471 : 1;
	1472 : 1;
	1473 : 1;
	1474 : 1;
	1475 : 1;
	1476 : 1;
	1477 : 1;
	1478 : 1;
	1479 : 1;
	1480 : 1;
	1481 : 1;
	1482 : 1;
	1483 : 1;
	1484 : 1;
	1485 : 1;
	1486 : 1;
	1487 : 1;
	1488 : 1;
	1489 : 1;
	1490 : 1;
	1491 : 1;
	1492 : 1;
	1493 : 1;
	1494 : 1;
	1495 : 1;
	1496 : 1;
	1497 : 1;
	1498 : 1;
	1499 : 1;
	1500 : 1;
	1501 : 1;
	1502 : 1;
	1503 : 1;
	1504 : 1;
	1505 : 1;
	1506 : 1;
	1507 : 1;
	1508 : 1;
	1509 : 1;
	1510 : 1;
	1511 : 1;
	1512 : 1;
	1513 : 1;
	1514 : 1;
	1515 : 1;
	1516 : 1;
	1517 : 1;
	1518 : 1;
	1519 : 1;
	1520 : 1;
	1521 : 1;
	1522 : 1;
	1523 : 1;
	1524 : 1;
	1525 : 1;
	1526 : 1;
	1527 : 1;
	1528 : 1;
	1529 : 1;
	1530 : 1;
	1531 : 1;
	1532 : 1;
	1533 : 1;
	1534 : 1;
	1535 : 1;
	1536 : 1;
	1537 : 1;
	1538 : 1;
	1539 : 1;
	1540 : 1;
	1541 : 1;
	1542 : 1;
	1543 : 1;
	1544 : 1;
	1545 : 1;
	1546 : 1;
	1547 : 1;
	1548 : 1;
	1549 : 1;
	1550 : 1;
	1551 : 1;
	1552 : 1;
	1553 : 1;
	1554 : 1;
	1555 : 1;
	1556 : 1;
	1557 : 1;
	1558 : 1;
	1559 : 1;
	1560 : 1;
	1561 : 1;
	1562 : 1;
	1563 : 1;
	1564 : 1;
	1565 : 1;
	1566 : 1;
	1567 : 1;
	1568 : 1;
	1569 : 1;
	1570 : 1;
	1571 : 1;
	1572 : 1;
	1573 : 1;
	1574 : 1;
	1575 : 1;
	1576 : 1;
	1577 : 1;
	1578 : 1;
	1579 : 1;
	1580 : 1;
	1581 : 1;
	1582 : 1;
	1583 : 1;
	1584 : 1;
	1585 : 1;
	1586 : 1;
	1587 : 1;
	1588 : 1;
	1589 : 1;
	1590 : 1;
	1591 : 1;
	1592 : 1;
	1593 : 1;
	1594 : 1;
	1595 : 1;
	1596 : 1;
	1597 : 1;
	1598 : 1;
	1599 : 1;
	1600 : 1;
	1601 : 1;
	1602 : 1;
	1603 : 1;
	1604 : 1;
	1605 : 1;
	1606 : 1;
	1607 : 1;
	1608 : 1;
	1609 : 1;
	1610 : 1;
	1611 : 1;
	1612 : 1;
	1613 : 1;
	1614 : 1;
	1615 : 1;
	1616 : 1;
	1617 : 1;
	1618 : 1;
	1619 : 1;
	1620 : 1;
	1621 : 1;
	1622 : 1;
	1623 : 1;
	1624 : 1;
	1625 : 1;
	1626 : 1;
	1627 : 1;
	1628 : 1;
	1629 : 1;
	1630 : 1;
	1631 : 1;
	1632 : 1;
	1633 : 1;
	1634 : 1;
	1635 : 1;
	1636 : 1;
	1637 : 1;
	1638 : 1;
	1639 : 1;
	1640 : 1;
	1641 : 1;
	1642 : 1;
	1643 : 1;
	1644 : 1;
	1645 : 1;
	1646 : 1;
	1647 : 1;
	1648 : 1;
	1649 : 1;
	1650 : 1;
	1651 : 1;
	1652 : 1;
	1653 : 1;
	1654 : 1;
	1655 : 1;
	1656 : 1;
	1657 : 1;
	1658 : 1;
	1659 : 1;
	1660 : 1;
	1661 : 1;
	1662 : 1;
	1663 : 1;
	1664 : 1;
	1665 : 1;
	1666 : 1;
	1667 : 1;
	1668 : 1;
	1669 : 1;
	1670 : 1;
	1671 : 1;
	1672 : 1;
	1673 : 1;
	1674 : 1;
	1675 : 1;
	1676 : 1;
	1677 : 1;
	1678 : 1;
	1679 : 1;
	1680 : 1;
	1681 : 1;
	1682 : 1;
	1683 : 1;
	1684 : 1;
	1685 : 1;
	1686 : 1;
	1687 : 1;
	1688 : 1;
	1689 : 1;
	1690 : 1;
	1691 : 1;
	1692 : 1;
	1693 : 1;
	1694 : 1;
	1695 : 1;
	1696 : 1;
	1697 : 1;
	1698 : 1;
	1699 : 1;
	1700 : 1;
	1701 : 1;
	1702 : 1;
	1703 : 1;
	1704 : 1;
	1705 : 1;
	1706 : 1;
	1707 : 1;
	1708 : 1;
	1709 : 1;
	1710 : 1;
	1711 : 1;
	1712 : 1;
	1713 : 1;
	1714 : 1;
	1715 : 1;
	1716 : 1;
	1717 : 1;
	1718 : 1;
	1719 : 1;
	1720 : 1;
	1721 : 1;
	1722 : 1;
	1723 : 1;
	1724 : 1;
	1725 : 1;
	1726 : 1;
	1727 : 1;
	1728 : 1;
	1729 : 1;
	1730 : 1;
	1731 : 1;
	1732 : 1;
	1733 : 1;
	1734 : 1;
	1735 : 1;
	1736 : 1;
	1737 : 1;
	1738 : 1;
	1739 : 1;
	1740 : 1;
	1741 : 1;
	1742 : 1;
	1743 : 1;
	1744 : 1;
	1745 : 1;
	1746 : 1;
	1747 : 1;
	1748 : 1;
	1749 : 1;
	1750 : 1;
	1751 : 1;
	1752 : 1;
	1753 : 1;
	1754 : 1;
	1755 : 1;
	1756 : 1;
	1757 : 1;
	1758 : 1;
	1759 : 1;
	1760 : 1;
	1761 : 1;
	1762 : 1;
	1763 : 1;
	1764 : 1;
	1765 : 1;
	1766 : 1;
	1767 : 1;
	1768 : 1;
	1769 : 1;
	1770 : 1;
	1771 : 1;
	1772 : 1;
	1773 : 1;
	1774 : 1;
	1775 : 1;
	1776 : 1;
	1777 : 1;
	1778 : 1;
	1779 : 1;
	1780 : 1;
	1781 : 1;
	1782 : 1;
	1783 : 1;
	1784 : 1;
	1785 : 1;
	1786 : 1;
	1787 : 1;
	1788 : 1;
	1789 : 1;
	1790 : 1;
	1791 : 1;
	1792 : 1;
	1793 : 1;
	1794 : 1;
	1795 : 1;
	1796 : 1;
	1797 : 1;
	1798 : 1;
	1799 : 1;
	1800 : 1;
	1801 : 1;
	1802 : 1;
	1803 : 1;
	1804 : 1;
	1805 : 1;
	1806 : 1;
	1807 : 1;
	1808 : 1;
	1809 : 1;
	1810 : 1;
	1811 : 1;
	1812 : 1;
	1813 : 1;
	1814 : 1;
	1815 : 1;
	1816 : 1;
	1817 : 1;
	1818 : 1;
	1819 : 1;
	1820 : 1;
	1821 : 1;
	1822 : 1;
	1823 : 1;
	1824 : 1;
	1825 : 1;
	1826 : 1;
	1827 : 1;
	1828 : 1;
	1829 : 1;
	1830 : 1;
	1831 : 1;
	1832 : 1;
	1833 : 1;
	1834 : 1;
	1835 : 1;
	1836 : 1;
	1837 : 1;
	1838 : 1;
	1839 : 1;
	1840 : 1;
	1841 : 1;
	1842 : 1;
	1843 : 1;
	1844 : 1;
	1845 : 1;
	1846 : 1;
	1847 : 1;
	1848 : 1;
	1849 : 1;
	1850 : 1;
	1851 : 1;
	1852 : 1;
	1853 : 1;
	1854 : 1;
	1855 : 1;
	1856 : 1;
	1857 : 1;
	1858 : 1;
	1859 : 1;
	1860 : 1;
	1861 : 1;
	1862 : 1;
	1863 : 1;
	1864 : 1;
	1865 : 1;
	1866 : 1;
	1867 : 1;
	1868 : 1;
	1869 : 1;
	1870 : 1;
	1871 : 1;
	1872 : 1;
	1873 : 1;
	1874 : 1;
	1875 : 1;
	1876 : 1;
	1877 : 1;
	1878 : 1;
	1879 : 1;
	1880 : 1;
	1881 : 1;
	1882 : 1;
	1883 : 1;
	1884 : 1;
	1885 : 1;
	1886 : 1;
	1887 : 1;
	1888 : 1;
	1889 : 1;
	1890 : 1;
	1891 : 1;
	1892 : 1;
	1893 : 1;
	1894 : 1;
	1895 : 1;
	1896 : 1;
	1897 : 1;
	1898 : 1;
	1899 : 1;
	1900 : 1;
	1901 : 1;
	1902 : 1;
	1903 : 1;
	1904 : 1;
	1905 : 1;
	1906 : 1;
	1907 : 1;
	1908 : 1;
	1909 : 1;
	1910 : 1;
	1911 : 1;
	1912 : 1;
	1913 : 1;
	1914 : 1;
	1915 : 1;
	1916 : 1;
	1917 : 1;
	1918 : 1;
	1919 : 1;
	1920 : 1;
	1921 : 1;
	1922 : 1;
	1923 : 1;
	1924 : 1;
	1925 : 1;
	1926 : 1;
	1927 : 1;
	1928 : 1;
	1929 : 1;
	1930 : 1;
	1931 : 1;
	1932 : 1;
	1933 : 1;
	1934 : 1;
	1935 : 1;
	1936 : 1;
	1937 : 1;
	1938 : 1;
	1939 : 1;
	1940 : 1;
	1941 : 1;
	1942 : 1;
	1943 : 1;
	1944 : 1;
	1945 : 1;
	1946 : 1;
	1947 : 1;
	1948 : 1;
	1949 : 1;
	1950 : 1;
	1951 : 1;
	1952 : 1;
	1953 : 1;
	1954 : 1;
	1955 : 1;
	1956 : 1;
	1957 : 1;
	1958 : 1;
	1959 : 1;
	1960 : 1;
	1961 : 1;
	1962 : 1;
	1963 : 1;
	1964 : 1;
	1965 : 1;
	1966 : 1;
	1967 : 1;
	1968 : 1;
	1969 : 1;
	1970 : 1;
	1971 : 1;
	1972 : 1;
	1973 : 1;
	1974 : 0;
	1975 : 1;
	1976 : 1;
	1977 : 1;
	1978 : 1;
	1979 : 1;
	1980 : 1;
	1981 : 1;
	1982 : 1;
	1983 : 1;
	1984 : 1;
	1985 : 1;
	1986 : 1;
	1987 : 1;
	1988 : 1;
	1989 : 1;
	1990 : 1;
	1991 : 1;
	1992 : 1;
	1993 : 1;
	1994 : 1;
	1995 : 1;
	1996 : 1;
	1997 : 1;
	1998 : 1;
	1999 : 1;
	2000 : 1;
	2001 : 1;
	2002 : 1;
	2003 : 1;
	2004 : 1;
	2005 : 1;
	2006 : 1;
	2007 : 1;
	2008 : 1;
	2009 : 1;
	2010 : 1;
	2011 : 1;
	2012 : 1;
	2013 : 1;
	2014 : 1;
	2015 : 1;
	2016 : 1;
	2017 : 1;
	2018 : 1;
	2019 : 1;
	2020 : 1;
	2021 : 1;
	2022 : 1;
	2023 : 1;
	2024 : 1;
	2025 : 1;
	2026 : 1;
	2027 : 1;
	2028 : 1;
	2029 : 1;
	2030 : 1;
	2031 : 1;
	2032 : 1;
	2033 : 1;
	2034 : 1;
	2035 : 1;
	2036 : 1;
	2037 : 1;
	2038 : 1;
	2039 : 1;
	2040 : 1;
	2041 : 1;
	2042 : 1;
	2043 : 1;
	2044 : 1;
	2045 : 1;
	2046 : 1;
	2047 : 1;
	2048 : 1;
	2049 : 1;
	2050 : 1;
	2051 : 1;
	2052 : 1;
	2053 : 1;
	2054 : 1;
	2055 : 1;
	2056 : 1;
	2057 : 1;
	2058 : 1;
	2059 : 1;
	2060 : 1;
	2061 : 1;
	2062 : 1;
	2063 : 1;
	2064 : 1;
	2065 : 1;
	2066 : 1;
	2067 : 1;
	2068 : 1;
	2069 : 1;
	2070 : 1;
	2071 : 1;
	2072 : 1;
	2073 : 1;
	2074 : 1;
	2075 : 1;
	2076 : 1;
	2077 : 1;
	2078 : 1;
	2079 : 1;
	2080 : 1;
	2081 : 1;
	2082 : 1;
	2083 : 1;
	2084 : 1;
	2085 : 1;
	2086 : 1;
	2087 : 1;
	2088 : 1;
	2089 : 1;
	2090 : 1;
	2091 : 1;
	2092 : 1;
	2093 : 1;
	2094 : 1;
	2095 : 1;
	2096 : 1;
	2097 : 1;
	2098 : 1;
	2099 : 1;
	2100 : 1;
	2101 : 1;
	2102 : 1;
	2103 : 1;
	2104 : 1;
	2105 : 1;
	2106 : 1;
	2107 : 1;
	2108 : 1;
	2109 : 1;
	2110 : 1;
	2111 : 1;
	2112 : 1;
	2113 : 1;
	2114 : 1;
	2115 : 1;
	2116 : 1;
	2117 : 1;
	2118 : 1;
	2119 : 1;
	2120 : 1;
	2121 : 1;
	2122 : 1;
	2123 : 1;
	2124 : 1;
	2125 : 1;
	2126 : 1;
	2127 : 1;
	2128 : 1;
	2129 : 1;
	2130 : 1;
	2131 : 1;
	2132 : 1;
	2133 : 1;
	2134 : 1;
	2135 : 1;
	2136 : 1;
	2137 : 1;
	2138 : 1;
	2139 : 1;
	2140 : 1;
	2141 : 1;
	2142 : 1;
	2143 : 1;
	2144 : 1;
	2145 : 1;
	2146 : 1;
	2147 : 1;
	2148 : 1;
	2149 : 1;
	2150 : 1;
	2151 : 1;
	2152 : 1;
	2153 : 1;
	2154 : 1;
	2155 : 1;
	2156 : 1;
	2157 : 1;
	2158 : 1;
	2159 : 1;
	2160 : 1;
	2161 : 1;
	2162 : 1;
	2163 : 1;
	2164 : 1;
	2165 : 1;
	2166 : 1;
	2167 : 1;
	2168 : 1;
	2169 : 1;
	2170 : 1;
	2171 : 1;
	2172 : 1;
	2173 : 1;
	2174 : 1;
	2175 : 1;
	2176 : 1;
	2177 : 1;
	2178 : 1;
	2179 : 1;
	2180 : 1;
	2181 : 1;
	2182 : 1;
	2183 : 1;
	2184 : 1;
	2185 : 1;
	2186 : 1;
	2187 : 1;
	2188 : 1;
	2189 : 1;
	2190 : 1;
	2191 : 1;
	2192 : 1;
	2193 : 1;
	2194 : 1;
	2195 : 1;
	2196 : 1;
	2197 : 1;
	2198 : 1;
	2199 : 1;
	2200 : 1;
	2201 : 1;
	2202 : 1;
	2203 : 1;
	2204 : 1;
	2205 : 1;
	2206 : 1;
	2207 : 1;
	2208 : 1;
	2209 : 1;
	2210 : 0;
	2211 : 1;
	2212 : 1;
	2213 : 0;
	2214 : 0;
	2215 : 1;
	2216 : 1;
	2217 : 1;
	2218 : 1;
	2219 : 1;
	2220 : 1;
	2221 : 1;
	2222 : 1;
	2223 : 1;
	2224 : 1;
	2225 : 1;
	2226 : 1;
	2227 : 1;
	2228 : 1;
	2229 : 1;
	2230 : 1;
	2231 : 1;
	2232 : 1;
	2233 : 1;
	2234 : 1;
	2235 : 1;
	2236 : 1;
	2237 : 1;
	2238 : 1;
	2239 : 1;
	2240 : 1;
	2241 : 1;
	2242 : 1;
	2243 : 1;
	2244 : 1;
	2245 : 1;
	2246 : 1;
	2247 : 1;
	2248 : 1;
	2249 : 1;
	2250 : 1;
	2251 : 1;
	2252 : 1;
	2253 : 1;
	2254 : 1;
	2255 : 1;
	2256 : 1;
	2257 : 1;
	2258 : 1;
	2259 : 1;
	2260 : 1;
	2261 : 1;
	2262 : 1;
	2263 : 1;
	2264 : 1;
	2265 : 1;
	2266 : 1;
	2267 : 1;
	2268 : 1;
	2269 : 1;
	2270 : 1;
	2271 : 1;
	2272 : 1;
	2273 : 1;
	2274 : 1;
	2275 : 1;
	2276 : 1;
	2277 : 1;
	2278 : 1;
	2279 : 1;
	2280 : 1;
	2281 : 1;
	2282 : 1;
	2283 : 1;
	2284 : 1;
	2285 : 1;
	2286 : 1;
	2287 : 1;
	2288 : 1;
	2289 : 1;
	2290 : 1;
	2291 : 1;
	2292 : 1;
	2293 : 1;
	2294 : 1;
	2295 : 1;
	2296 : 1;
	2297 : 1;
	2298 : 1;
	2299 : 1;
	2300 : 1;
	2301 : 1;
	2302 : 1;
	2303 : 1;
	2304 : 1;
	2305 : 1;
	2306 : 1;
	2307 : 1;
	2308 : 1;
	2309 : 1;
	2310 : 1;
	2311 : 1;
	2312 : 1;
	2313 : 1;
	2314 : 1;
	2315 : 1;
	2316 : 1;
	2317 : 1;
	2318 : 1;
	2319 : 1;
	2320 : 1;
	2321 : 1;
	2322 : 1;
	2323 : 1;
	2324 : 1;
	2325 : 1;
	2326 : 1;
	2327 : 1;
	2328 : 1;
	2329 : 1;
	2330 : 1;
	2331 : 1;
	2332 : 1;
	2333 : 1;
	2334 : 1;
	2335 : 1;
	2336 : 1;
	2337 : 1;
	2338 : 1;
	2339 : 1;
	2340 : 1;
	2341 : 1;
	2342 : 1;
	2343 : 1;
	2344 : 1;
	2345 : 1;
	2346 : 1;
	2347 : 1;
	2348 : 1;
	2349 : 1;
	2350 : 1;
	2351 : 1;
	2352 : 1;
	2353 : 1;
	2354 : 1;
	2355 : 1;
	2356 : 1;
	2357 : 1;
	2358 : 1;
	2359 : 1;
	2360 : 1;
	2361 : 1;
	2362 : 1;
	2363 : 1;
	2364 : 1;
	2365 : 1;
	2366 : 1;
	2367 : 1;
	2368 : 1;
	2369 : 1;
	2370 : 1;
	2371 : 1;
	2372 : 1;
	2373 : 1;
	2374 : 1;
	2375 : 1;
	2376 : 1;
	2377 : 1;
	2378 : 1;
	2379 : 1;
	2380 : 1;
	2381 : 1;
	2382 : 1;
	2383 : 1;
	2384 : 1;
	2385 : 1;
	2386 : 1;
	2387 : 1;
	2388 : 1;
	2389 : 1;
	2390 : 1;
	2391 : 1;
	2392 : 1;
	2393 : 1;
	2394 : 1;
	2395 : 1;
	2396 : 1;
	2397 : 1;
	2398 : 1;
	2399 : 1;
	2400 : 1;
	2401 : 1;
	2402 : 1;
	2403 : 1;
	2404 : 1;
	2405 : 1;
	2406 : 1;
	2407 : 1;
	2408 : 1;
	2409 : 1;
	2410 : 1;
	2411 : 1;
	2412 : 1;
	2413 : 1;
	2414 : 1;
	2415 : 1;
	2416 : 1;
	2417 : 1;
	2418 : 1;
	2419 : 1;
	2420 : 1;
	2421 : 1;
	2422 : 1;
	2423 : 1;
	2424 : 1;
	2425 : 1;
	2426 : 1;
	2427 : 1;
	2428 : 1;
	2429 : 1;
	2430 : 1;
	2431 : 1;
	2432 : 1;
	2433 : 1;
	2434 : 1;
	2435 : 1;
	2436 : 1;
	2437 : 1;
	2438 : 1;
	2439 : 1;
	2440 : 1;
	2441 : 1;
	2442 : 1;
	2443 : 1;
	2444 : 1;
	2445 : 1;
	2446 : 1;
	2447 : 1;
	2448 : 1;
	2449 : 1;
	2450 : 0;
	2451 : 1;
	2452 : 1;
	2453 : 0;
	2454 : 0;
	2455 : 1;
	2456 : 1;
	2457 : 1;
	2458 : 1;
	2459 : 1;
	2460 : 1;
	2461 : 1;
	2462 : 1;
	2463 : 1;
	2464 : 1;
	2465 : 1;
	2466 : 1;
	2467 : 1;
	2468 : 1;
	2469 : 1;
	2470 : 1;
	2471 : 1;
	2472 : 1;
	2473 : 1;
	2474 : 1;
	2475 : 1;
	2476 : 1;
	2477 : 1;
	2478 : 1;
	2479 : 1;
	2480 : 1;
	2481 : 1;
	2482 : 1;
	2483 : 1;
	2484 : 1;
	2485 : 1;
	2486 : 1;
	2487 : 1;
	2488 : 1;
	2489 : 1;
	2490 : 1;
	2491 : 1;
	2492 : 1;
	2493 : 1;
	2494 : 1;
	2495 : 1;
	2496 : 1;
	2497 : 1;
	2498 : 1;
	2499 : 1;
	2500 : 1;
	2501 : 1;
	2502 : 1;
	2503 : 1;
	2504 : 1;
	2505 : 1;
	2506 : 1;
	2507 : 1;
	2508 : 1;
	2509 : 1;
	2510 : 1;
	2511 : 1;
	2512 : 1;
	2513 : 1;
	2514 : 1;
	2515 : 1;
	2516 : 1;
	2517 : 1;
	2518 : 1;
	2519 : 1;
	2520 : 1;
	2521 : 1;
	2522 : 1;
	2523 : 1;
	2524 : 1;
	2525 : 1;
	2526 : 1;
	2527 : 1;
	2528 : 1;
	2529 : 1;
	2530 : 1;
	2531 : 1;
	2532 : 1;
	2533 : 1;
	2534 : 1;
	2535 : 1;
	2536 : 1;
	2537 : 1;
	2538 : 1;
	2539 : 1;
	2540 : 1;
	2541 : 1;
	2542 : 1;
	2543 : 1;
	2544 : 1;
	2545 : 1;
	2546 : 1;
	2547 : 1;
	2548 : 1;
	2549 : 1;
	2550 : 1;
	2551 : 1;
	2552 : 1;
	2553 : 1;
	2554 : 1;
	2555 : 1;
	2556 : 1;
	2557 : 1;
	2558 : 1;
	2559 : 1;
	2560 : 1;
	2561 : 1;
	2562 : 1;
	2563 : 1;
	2564 : 1;
	2565 : 1;
	2566 : 1;
	2567 : 1;
	2568 : 1;
	2569 : 1;
	2570 : 1;
	2571 : 1;
	2572 : 1;
	2573 : 1;
	2574 : 1;
	2575 : 1;
	2576 : 1;
	2577 : 1;
	2578 : 1;
	2579 : 1;
	2580 : 1;
	2581 : 1;
	2582 : 1;
	2583 : 1;
	2584 : 1;
	2585 : 1;
	2586 : 1;
	2587 : 1;
	2588 : 1;
	2589 : 1;
	2590 : 1;
	2591 : 1;
	2592 : 1;
	2593 : 1;
	2594 : 1;
	2595 : 1;
	2596 : 1;
	2597 : 1;
	2598 : 1;
	2599 : 1;
	2600 : 1;
	2601 : 1;
	2602 : 1;
	2603 : 1;
	2604 : 1;
	2605 : 1;
	2606 : 1;
	2607 : 1;
	2608 : 1;
	2609 : 1;
	2610 : 1;
	2611 : 1;
	2612 : 1;
	2613 : 1;
	2614 : 1;
	2615 : 1;
	2616 : 1;
	2617 : 1;
	2618 : 1;
	2619 : 1;
	2620 : 1;
	2621 : 1;
	2622 : 1;
	2623 : 1;
	2624 : 1;
	2625 : 1;
	2626 : 1;
	2627 : 1;
	2628 : 1;
	2629 : 1;
	2630 : 1;
	2631 : 1;
	2632 : 1;
	2633 : 1;
	2634 : 1;
	2635 : 1;
	2636 : 1;
	2637 : 1;
	2638 : 1;
	2639 : 1;
	2640 : 1;
	2641 : 1;
	2642 : 1;
	2643 : 1;
	2644 : 1;
	2645 : 1;
	2646 : 1;
	2647 : 1;
	2648 : 1;
	2649 : 1;
	2650 : 1;
	2651 : 1;
	2652 : 1;
	2653 : 1;
	2654 : 1;
	2655 : 1;
	2656 : 1;
	2657 : 1;
	2658 : 1;
	2659 : 1;
	2660 : 1;
	2661 : 1;
	2662 : 1;
	2663 : 1;
	2664 : 1;
	2665 : 1;
	2666 : 1;
	2667 : 1;
	2668 : 1;
	2669 : 1;
	2670 : 1;
	2671 : 1;
	2672 : 1;
	2673 : 1;
	2674 : 1;
	2675 : 1;
	2676 : 1;
	2677 : 1;
	2678 : 1;
	2679 : 1;
	2680 : 1;
	2681 : 1;
	2682 : 1;
	2683 : 1;
	2684 : 1;
	2685 : 1;
	2686 : 1;
	2687 : 1;
	2688 : 1;
	2689 : 1;
	2690 : 0;
	2691 : 0;
	2692 : 1;
	2693 : 0;
	2694 : 0;
	2695 : 1;
	2696 : 1;
	2697 : 1;
	2698 : 1;
	2699 : 1;
	2700 : 1;
	2701 : 1;
	2702 : 1;
	2703 : 1;
	2704 : 1;
	2705 : 1;
	2706 : 1;
	2707 : 1;
	2708 : 1;
	2709 : 1;
	2710 : 1;
	2711 : 1;
	2712 : 1;
	2713 : 1;
	2714 : 1;
	2715 : 1;
	2716 : 1;
	2717 : 1;
	2718 : 1;
	2719 : 1;
	2720 : 1;
	2721 : 1;
	2722 : 1;
	2723 : 1;
	2724 : 1;
	2725 : 1;
	2726 : 1;
	2727 : 1;
	2728 : 1;
	2729 : 1;
	2730 : 1;
	2731 : 1;
	2732 : 1;
	2733 : 1;
	2734 : 1;
	2735 : 1;
	2736 : 1;
	2737 : 1;
	2738 : 1;
	2739 : 1;
	2740 : 1;
	2741 : 1;
	2742 : 0;
	2743 : 1;
	2744 : 1;
	2745 : 1;
	2746 : 1;
	2747 : 1;
	2748 : 1;
	2749 : 1;
	2750 : 1;
	2751 : 1;
	2752 : 1;
	2753 : 1;
	2754 : 1;
	2755 : 1;
	2756 : 1;
	2757 : 1;
	2758 : 1;
	2759 : 1;
	2760 : 1;
	2761 : 1;
	2762 : 1;
	2763 : 1;
	2764 : 1;
	2765 : 1;
	2766 : 1;
	2767 : 1;
	2768 : 1;
	2769 : 1;
	2770 : 1;
	2771 : 1;
	2772 : 1;
	2773 : 1;
	2774 : 1;
	2775 : 1;
	2776 : 1;
	2777 : 1;
	2778 : 1;
	2779 : 1;
	2780 : 1;
	2781 : 1;
	2782 : 1;
	2783 : 1;
	2784 : 1;
	2785 : 1;
	2786 : 1;
	2787 : 1;
	2788 : 1;
	2789 : 1;
	2790 : 1;
	2791 : 1;
	2792 : 1;
	2793 : 1;
	2794 : 1;
	2795 : 1;
	2796 : 1;
	2797 : 1;
	2798 : 1;
	2799 : 1;
	2800 : 1;
	2801 : 1;
	2802 : 1;
	2803 : 1;
	2804 : 1;
	2805 : 1;
	2806 : 1;
	2807 : 1;
	2808 : 1;
	2809 : 1;
	2810 : 1;
	2811 : 1;
	2812 : 1;
	2813 : 1;
	2814 : 1;
	2815 : 1;
	2816 : 1;
	2817 : 1;
	2818 : 1;
	2819 : 1;
	2820 : 1;
	2821 : 1;
	2822 : 1;
	2823 : 1;
	2824 : 1;
	2825 : 1;
	2826 : 1;
	2827 : 1;
	2828 : 1;
	2829 : 1;
	2830 : 1;
	2831 : 1;
	2832 : 1;
	2833 : 1;
	2834 : 1;
	2835 : 1;
	2836 : 1;
	2837 : 1;
	2838 : 1;
	2839 : 1;
	2840 : 1;
	2841 : 1;
	2842 : 1;
	2843 : 1;
	2844 : 1;
	2845 : 1;
	2846 : 0;
	2847 : 0;
	2848 : 0;
	2849 : 1;
	2850 : 1;
	2851 : 1;
	2852 : 1;
	2853 : 0;
	2854 : 0;
	2855 : 1;
	2856 : 1;
	2857 : 1;
	2858 : 0;
	2859 : 0;
	2860 : 0;
	2861 : 0;
	2862 : 1;
	2863 : 1;
	2864 : 1;
	2865 : 1;
	2866 : 1;
	2867 : 1;
	2868 : 1;
	2869 : 1;
	2870 : 1;
	2871 : 1;
	2872 : 1;
	2873 : 1;
	2874 : 1;
	2875 : 1;
	2876 : 1;
	2877 : 1;
	2878 : 1;
	2879 : 1;
	2880 : 1;
	2881 : 1;
	2882 : 1;
	2883 : 1;
	2884 : 1;
	2885 : 1;
	2886 : 1;
	2887 : 1;
	2888 : 1;
	2889 : 1;
	2890 : 1;
	2891 : 1;
	2892 : 1;
	2893 : 1;
	2894 : 1;
	2895 : 1;
	2896 : 1;
	2897 : 1;
	2898 : 1;
	2899 : 1;
	2900 : 1;
	2901 : 1;
	2902 : 1;
	2903 : 1;
	2904 : 1;
	2905 : 1;
	2906 : 1;
	2907 : 1;
	2908 : 1;
	2909 : 1;
	2910 : 1;
	2911 : 1;
	2912 : 1;
	2913 : 1;
	2914 : 1;
	2915 : 1;
	2916 : 1;
	2917 : 1;
	2918 : 1;
	2919 : 1;
	2920 : 1;
	2921 : 1;
	2922 : 1;
	2923 : 1;
	2924 : 1;
	2925 : 1;
	2926 : 1;
	2927 : 1;
	2928 : 1;
	2929 : 1;
	2930 : 0;
	2931 : 0;
	2932 : 1;
	2933 : 0;
	2934 : 0;
	2935 : 1;
	2936 : 1;
	2937 : 1;
	2938 : 1;
	2939 : 1;
	2940 : 1;
	2941 : 1;
	2942 : 1;
	2943 : 1;
	2944 : 1;
	2945 : 1;
	2946 : 1;
	2947 : 1;
	2948 : 1;
	2949 : 1;
	2950 : 1;
	2951 : 1;
	2952 : 1;
	2953 : 1;
	2954 : 1;
	2955 : 1;
	2956 : 1;
	2957 : 1;
	2958 : 1;
	2959 : 1;
	2960 : 1;
	2961 : 1;
	2962 : 1;
	2963 : 1;
	2964 : 1;
	2965 : 1;
	2966 : 1;
	2967 : 1;
	2968 : 1;
	2969 : 1;
	2970 : 1;
	2971 : 1;
	2972 : 1;
	2973 : 1;
	2974 : 1;
	2975 : 1;
	2976 : 1;
	2977 : 1;
	2978 : 1;
	2979 : 1;
	2980 : 1;
	2981 : 1;
	2982 : 0;
	2983 : 1;
	2984 : 1;
	2985 : 1;
	2986 : 1;
	2987 : 1;
	2988 : 1;
	2989 : 1;
	2990 : 1;
	2991 : 1;
	2992 : 1;
	2993 : 1;
	2994 : 1;
	2995 : 1;
	2996 : 1;
	2997 : 1;
	2998 : 1;
	2999 : 1;
	3000 : 1;
	3001 : 1;
	3002 : 1;
	3003 : 1;
	3004 : 1;
	3005 : 1;
	3006 : 1;
	3007 : 1;
	3008 : 1;
	3009 : 1;
	3010 : 1;
	3011 : 1;
	3012 : 1;
	3013 : 1;
	3014 : 1;
	3015 : 1;
	3016 : 1;
	3017 : 1;
	3018 : 1;
	3019 : 1;
	3020 : 1;
	3021 : 1;
	3022 : 1;
	3023 : 1;
	3024 : 1;
	3025 : 1;
	3026 : 1;
	3027 : 1;
	3028 : 1;
	3029 : 1;
	3030 : 1;
	3031 : 1;
	3032 : 1;
	3033 : 1;
	3034 : 1;
	3035 : 1;
	3036 : 1;
	3037 : 1;
	3038 : 1;
	3039 : 1;
	3040 : 1;
	3041 : 1;
	3042 : 1;
	3043 : 1;
	3044 : 1;
	3045 : 1;
	3046 : 1;
	3047 : 1;
	3048 : 1;
	3049 : 1;
	3050 : 1;
	3051 : 1;
	3052 : 1;
	3053 : 1;
	3054 : 1;
	3055 : 1;
	3056 : 1;
	3057 : 1;
	3058 : 1;
	3059 : 1;
	3060 : 1;
	3061 : 1;
	3062 : 1;
	3063 : 1;
	3064 : 1;
	3065 : 1;
	3066 : 1;
	3067 : 1;
	3068 : 1;
	3069 : 1;
	3070 : 1;
	3071 : 1;
	3072 : 1;
	3073 : 1;
	3074 : 1;
	3075 : 1;
	3076 : 1;
	3077 : 1;
	3078 : 1;
	3079 : 1;
	3080 : 1;
	3081 : 1;
	3082 : 1;
	3083 : 1;
	3084 : 1;
	3085 : 1;
	3086 : 0;
	3087 : 0;
	3088 : 0;
	3089 : 0;
	3090 : 1;
	3091 : 1;
	3092 : 0;
	3093 : 0;
	3094 : 0;
	3095 : 0;
	3096 : 1;
	3097 : 0;
	3098 : 0;
	3099 : 0;
	3100 : 0;
	3101 : 0;
	3102 : 0;
	3103 : 1;
	3104 : 1;
	3105 : 1;
	3106 : 1;
	3107 : 1;
	3108 : 1;
	3109 : 1;
	3110 : 1;
	3111 : 1;
	3112 : 1;
	3113 : 1;
	3114 : 1;
	3115 : 1;
	3116 : 1;
	3117 : 1;
	3118 : 1;
	3119 : 1;
	3120 : 1;
	3121 : 1;
	3122 : 1;
	3123 : 1;
	3124 : 1;
	3125 : 1;
	3126 : 1;
	3127 : 1;
	3128 : 1;
	3129 : 1;
	3130 : 1;
	3131 : 1;
	3132 : 1;
	3133 : 1;
	3134 : 0;
	3135 : 0;
	3136 : 0;
	3137 : 0;
	3138 : 0;
	3139 : 0;
	3140 : 1;
	3141 : 1;
	3142 : 1;
	3143 : 1;
	3144 : 1;
	3145 : 1;
	3146 : 1;
	3147 : 1;
	3148 : 1;
	3149 : 1;
	3150 : 1;
	3151 : 1;
	3152 : 1;
	3153 : 1;
	3154 : 1;
	3155 : 0;
	3156 : 0;
	3157 : 1;
	3158 : 1;
	3159 : 1;
	3160 : 1;
	3161 : 1;
	3162 : 1;
	3163 : 1;
	3164 : 1;
	3165 : 1;
	3166 : 1;
	3167 : 1;
	3168 : 1;
	3169 : 1;
	3170 : 1;
	3171 : 1;
	3172 : 1;
	3173 : 1;
	3174 : 1;
	3175 : 1;
	3176 : 1;
	3177 : 0;
	3178 : 0;
	3179 : 0;
	3180 : 0;
	3181 : 1;
	3182 : 1;
	3183 : 1;
	3184 : 1;
	3185 : 1;
	3186 : 1;
	3187 : 1;
	3188 : 1;
	3189 : 1;
	3190 : 1;
	3191 : 1;
	3192 : 1;
	3193 : 1;
	3194 : 1;
	3195 : 1;
	3196 : 1;
	3197 : 1;
	3198 : 1;
	3199 : 1;
	3200 : 1;
	3201 : 1;
	3202 : 1;
	3203 : 1;
	3204 : 1;
	3205 : 1;
	3206 : 1;
	3207 : 1;
	3208 : 1;
	3209 : 1;
	3210 : 1;
	3211 : 1;
	3212 : 1;
	3213 : 1;
	3214 : 1;
	3215 : 1;
	3216 : 1;
	3217 : 1;
	3218 : 1;
	3219 : 1;
	3220 : 1;
	3221 : 1;
	3222 : 0;
	3223 : 1;
	3224 : 1;
	3225 : 1;
	3226 : 0;
	3227 : 1;
	3228 : 1;
	3229 : 1;
	3230 : 0;
	3231 : 1;
	3232 : 1;
	3233 : 1;
	3234 : 1;
	3235 : 1;
	3236 : 1;
	3237 : 1;
	3238 : 1;
	3239 : 1;
	3240 : 1;
	3241 : 1;
	3242 : 1;
	3243 : 1;
	3244 : 1;
	3245 : 1;
	3246 : 1;
	3247 : 1;
	3248 : 1;
	3249 : 1;
	3250 : 1;
	3251 : 1;
	3252 : 1;
	3253 : 1;
	3254 : 1;
	3255 : 1;
	3256 : 1;
	3257 : 1;
	3258 : 1;
	3259 : 1;
	3260 : 1;
	3261 : 1;
	3262 : 1;
	3263 : 1;
	3264 : 1;
	3265 : 1;
	3266 : 1;
	3267 : 1;
	3268 : 1;
	3269 : 1;
	3270 : 1;
	3271 : 1;
	3272 : 1;
	3273 : 1;
	3274 : 1;
	3275 : 1;
	3276 : 1;
	3277 : 1;
	3278 : 1;
	3279 : 1;
	3280 : 1;
	3281 : 0;
	3282 : 0;
	3283 : 0;
	3284 : 0;
	3285 : 1;
	3286 : 1;
	3287 : 1;
	3288 : 1;
	3289 : 1;
	3290 : 1;
	3291 : 1;
	3292 : 1;
	3293 : 1;
	3294 : 1;
	3295 : 0;
	3296 : 1;
	3297 : 1;
	3298 : 1;
	3299 : 1;
	3300 : 1;
	3301 : 1;
	3302 : 1;
	3303 : 1;
	3304 : 0;
	3305 : 0;
	3306 : 0;
	3307 : 0;
	3308 : 0;
	3309 : 1;
	3310 : 1;
	3311 : 0;
	3312 : 0;
	3313 : 0;
	3314 : 0;
	3315 : 1;
	3316 : 0;
	3317 : 0;
	3318 : 0;
	3319 : 0;
	3320 : 0;
	3321 : 0;
	3322 : 1;
	3323 : 1;
	3324 : 1;
	3325 : 0;
	3326 : 1;
	3327 : 1;
	3328 : 1;
	3329 : 0;
	3330 : 1;
	3331 : 0;
	3332 : 1;
	3333 : 1;
	3334 : 1;
	3335 : 0;
	3336 : 0;
	3337 : 0;
	3338 : 0;
	3339 : 1;
	3340 : 1;
	3341 : 1;
	3342 : 1;
	3343 : 1;
	3344 : 1;
	3345 : 1;
	3346 : 1;
	3347 : 1;
	3348 : 1;
	3349 : 1;
	3350 : 1;
	3351 : 1;
	3352 : 1;
	3353 : 1;
	3354 : 1;
	3355 : 1;
	3356 : 1;
	3357 : 1;
	3358 : 1;
	3359 : 1;
	3360 : 1;
	3361 : 1;
	3362 : 1;
	3363 : 1;
	3364 : 1;
	3365 : 1;
	3366 : 1;
	3367 : 1;
	3368 : 1;
	3369 : 1;
	3370 : 1;
	3371 : 1;
	3372 : 1;
	3373 : 1;
	3374 : 1;
	3375 : 1;
	3376 : 1;
	3377 : 1;
	3378 : 0;
	3379 : 1;
	3380 : 1;
	3381 : 1;
	3382 : 1;
	3383 : 1;
	3384 : 1;
	3385 : 1;
	3386 : 1;
	3387 : 1;
	3388 : 1;
	3389 : 1;
	3390 : 1;
	3391 : 1;
	3392 : 1;
	3393 : 1;
	3394 : 0;
	3395 : 1;
	3396 : 1;
	3397 : 1;
	3398 : 1;
	3399 : 1;
	3400 : 1;
	3401 : 1;
	3402 : 1;
	3403 : 1;
	3404 : 0;
	3405 : 0;
	3406 : 0;
	3407 : 1;
	3408 : 1;
	3409 : 1;
	3410 : 1;
	3411 : 1;
	3412 : 1;
	3413 : 1;
	3414 : 1;
	3415 : 1;
	3416 : 0;
	3417 : 1;
	3418 : 1;
	3419 : 1;
	3420 : 0;
	3421 : 1;
	3422 : 1;
	3423 : 1;
	3424 : 1;
	3425 : 1;
	3426 : 1;
	3427 : 1;
	3428 : 1;
	3429 : 1;
	3430 : 1;
	3431 : 1;
	3432 : 1;
	3433 : 1;
	3434 : 1;
	3435 : 1;
	3436 : 1;
	3437 : 1;
	3438 : 1;
	3439 : 1;
	3440 : 1;
	3441 : 1;
	3442 : 1;
	3443 : 1;
	3444 : 1;
	3445 : 1;
	3446 : 1;
	3447 : 1;
	3448 : 1;
	3449 : 1;
	3450 : 1;
	3451 : 1;
	3452 : 0;
	3453 : 0;
	3454 : 1;
	3455 : 1;
	3456 : 1;
	3457 : 1;
	3458 : 1;
	3459 : 1;
	3460 : 1;
	3461 : 1;
	3462 : 0;
	3463 : 1;
	3464 : 1;
	3465 : 1;
	3466 : 0;
	3467 : 1;
	3468 : 1;
	3469 : 1;
	3470 : 0;
	3471 : 1;
	3472 : 1;
	3473 : 1;
	3474 : 1;
	3475 : 1;
	3476 : 1;
	3477 : 1;
	3478 : 1;
	3479 : 1;
	3480 : 1;
	3481 : 1;
	3482 : 1;
	3483 : 1;
	3484 : 1;
	3485 : 1;
	3486 : 1;
	3487 : 1;
	3488 : 1;
	3489 : 1;
	3490 : 1;
	3491 : 1;
	3492 : 1;
	3493 : 1;
	3494 : 1;
	3495 : 1;
	3496 : 1;
	3497 : 1;
	3498 : 1;
	3499 : 1;
	3500 : 0;
	3501 : 1;
	3502 : 1;
	3503 : 1;
	3504 : 1;
	3505 : 1;
	3506 : 1;
	3507 : 1;
	3508 : 1;
	3509 : 1;
	3510 : 1;
	3511 : 1;
	3512 : 1;
	3513 : 1;
	3514 : 1;
	3515 : 1;
	3516 : 1;
	3517 : 1;
	3518 : 1;
	3519 : 1;
	3520 : 0;
	3521 : 1;
	3522 : 1;
	3523 : 1;
	3524 : 0;
	3525 : 0;
	3526 : 1;
	3527 : 1;
	3528 : 0;
	3529 : 0;
	3530 : 1;
	3531 : 1;
	3532 : 1;
	3533 : 1;
	3534 : 1;
	3535 : 1;
	3536 : 1;
	3537 : 1;
	3538 : 1;
	3539 : 1;
	3540 : 1;
	3541 : 1;
	3542 : 1;
	3543 : 1;
	3544 : 0;
	3545 : 1;
	3546 : 1;
	3547 : 1;
	3548 : 1;
	3549 : 1;
	3550 : 0;
	3551 : 1;
	3552 : 1;
	3553 : 1;
	3554 : 1;
	3555 : 1;
	3556 : 0;
	3557 : 0;
	3558 : 1;
	3559 : 1;
	3560 : 1;
	3561 : 1;
	3562 : 1;
	3563 : 1;
	3564 : 1;
	3565 : 1;
	3566 : 1;
	3567 : 1;
	3568 : 1;
	3569 : 0;
	3570 : 1;
	3571 : 0;
	3572 : 1;
	3573 : 1;
	3574 : 1;
	3575 : 0;
	3576 : 0;
	3577 : 0;
	3578 : 0;
	3579 : 1;
	3580 : 1;
	3581 : 1;
	3582 : 1;
	3583 : 1;
	3584 : 1;
	3585 : 1;
	3586 : 1;
	3587 : 1;
	3588 : 1;
	3589 : 1;
	3590 : 1;
	3591 : 1;
	3592 : 1;
	3593 : 1;
	3594 : 1;
	3595 : 1;
	3596 : 1;
	3597 : 1;
	3598 : 1;
	3599 : 1;
	3600 : 1;
	3601 : 1;
	3602 : 1;
	3603 : 1;
	3604 : 1;
	3605 : 1;
	3606 : 1;
	3607 : 1;
	3608 : 1;
	3609 : 1;
	3610 : 1;
	3611 : 1;
	3612 : 1;
	3613 : 1;
	3614 : 1;
	3615 : 1;
	3616 : 1;
	3617 : 0;
	3618 : 1;
	3619 : 1;
	3620 : 1;
	3621 : 1;
	3622 : 1;
	3623 : 1;
	3624 : 1;
	3625 : 1;
	3626 : 1;
	3627 : 1;
	3628 : 1;
	3629 : 1;
	3630 : 1;
	3631 : 1;
	3632 : 1;
	3633 : 1;
	3634 : 0;
	3635 : 1;
	3636 : 1;
	3637 : 1;
	3638 : 1;
	3639 : 1;
	3640 : 1;
	3641 : 1;
	3642 : 1;
	3643 : 1;
	3644 : 1;
	3645 : 0;
	3646 : 1;
	3647 : 1;
	3648 : 1;
	3649 : 1;
	3650 : 1;
	3651 : 1;
	3652 : 1;
	3653 : 1;
	3654 : 1;
	3655 : 1;
	3656 : 0;
	3657 : 1;
	3658 : 1;
	3659 : 1;
	3660 : 1;
	3661 : 1;
	3662 : 1;
	3663 : 1;
	3664 : 1;
	3665 : 1;
	3666 : 1;
	3667 : 1;
	3668 : 1;
	3669 : 1;
	3670 : 1;
	3671 : 1;
	3672 : 1;
	3673 : 1;
	3674 : 1;
	3675 : 1;
	3676 : 1;
	3677 : 1;
	3678 : 1;
	3679 : 1;
	3680 : 1;
	3681 : 1;
	3682 : 1;
	3683 : 1;
	3684 : 1;
	3685 : 1;
	3686 : 1;
	3687 : 1;
	3688 : 1;
	3689 : 1;
	3690 : 1;
	3691 : 1;
	3692 : 0;
	3693 : 0;
	3694 : 1;
	3695 : 1;
	3696 : 1;
	3697 : 1;
	3698 : 1;
	3699 : 1;
	3700 : 1;
	3701 : 1;
	3702 : 0;
	3703 : 1;
	3704 : 1;
	3705 : 1;
	3706 : 1;
	3707 : 0;
	3708 : 1;
	3709 : 0;
	3710 : 1;
	3711 : 1;
	3712 : 1;
	3713 : 1;
	3714 : 1;
	3715 : 1;
	3716 : 1;
	3717 : 1;
	3718 : 1;
	3719 : 1;
	3720 : 1;
	3721 : 1;
	3722 : 1;
	3723 : 1;
	3724 : 1;
	3725 : 1;
	3726 : 1;
	3727 : 1;
	3728 : 1;
	3729 : 1;
	3730 : 1;
	3731 : 1;
	3732 : 1;
	3733 : 1;
	3734 : 1;
	3735 : 1;
	3736 : 1;
	3737 : 1;
	3738 : 1;
	3739 : 1;
	3740 : 0;
	3741 : 0;
	3742 : 1;
	3743 : 1;
	3744 : 1;
	3745 : 1;
	3746 : 1;
	3747 : 1;
	3748 : 1;
	3749 : 1;
	3750 : 1;
	3751 : 1;
	3752 : 1;
	3753 : 1;
	3754 : 1;
	3755 : 1;
	3756 : 1;
	3757 : 1;
	3758 : 1;
	3759 : 1;
	3760 : 0;
	3761 : 1;
	3762 : 1;
	3763 : 1;
	3764 : 0;
	3765 : 0;
	3766 : 1;
	3767 : 1;
	3768 : 0;
	3769 : 0;
	3770 : 1;
	3771 : 1;
	3772 : 1;
	3773 : 1;
	3774 : 1;
	3775 : 1;
	3776 : 1;
	3777 : 1;
	3778 : 1;
	3779 : 1;
	3780 : 1;
	3781 : 1;
	3782 : 1;
	3783 : 1;
	3784 : 0;
	3785 : 1;
	3786 : 1;
	3787 : 1;
	3788 : 1;
	3789 : 1;
	3790 : 0;
	3791 : 1;
	3792 : 1;
	3793 : 1;
	3794 : 1;
	3795 : 1;
	3796 : 0;
	3797 : 0;
	3798 : 1;
	3799 : 1;
	3800 : 1;
	3801 : 1;
	3802 : 1;
	3803 : 1;
	3804 : 1;
	3805 : 1;
	3806 : 1;
	3807 : 1;
	3808 : 1;
	3809 : 0;
	3810 : 1;
	3811 : 0;
	3812 : 0;
	3813 : 1;
	3814 : 1;
	3815 : 0;
	3816 : 1;
	3817 : 0;
	3818 : 0;
	3819 : 1;
	3820 : 1;
	3821 : 1;
	3822 : 1;
	3823 : 1;
	3824 : 1;
	3825 : 1;
	3826 : 1;
	3827 : 1;
	3828 : 1;
	3829 : 1;
	3830 : 1;
	3831 : 1;
	3832 : 1;
	3833 : 1;
	3834 : 1;
	3835 : 1;
	3836 : 1;
	3837 : 1;
	3838 : 1;
	3839 : 1;
	3840 : 1;
	3841 : 1;
	3842 : 1;
	3843 : 1;
	3844 : 1;
	3845 : 1;
	3846 : 1;
	3847 : 1;
	3848 : 1;
	3849 : 1;
	3850 : 1;
	3851 : 1;
	3852 : 1;
	3853 : 1;
	3854 : 1;
	3855 : 1;
	3856 : 0;
	3857 : 0;
	3858 : 1;
	3859 : 1;
	3860 : 0;
	3861 : 0;
	3862 : 1;
	3863 : 0;
	3864 : 0;
	3865 : 1;
	3866 : 1;
	3867 : 0;
	3868 : 0;
	3869 : 0;
	3870 : 0;
	3871 : 1;
	3872 : 1;
	3873 : 0;
	3874 : 0;
	3875 : 0;
	3876 : 0;
	3877 : 1;
	3878 : 0;
	3879 : 1;
	3880 : 1;
	3881 : 0;
	3882 : 0;
	3883 : 1;
	3884 : 1;
	3885 : 1;
	3886 : 1;
	3887 : 1;
	3888 : 1;
	3889 : 1;
	3890 : 1;
	3891 : 1;
	3892 : 1;
	3893 : 1;
	3894 : 1;
	3895 : 1;
	3896 : 0;
	3897 : 1;
	3898 : 1;
	3899 : 1;
	3900 : 1;
	3901 : 1;
	3902 : 1;
	3903 : 0;
	3904 : 0;
	3905 : 0;
	3906 : 0;
	3907 : 1;
	3908 : 0;
	3909 : 0;
	3910 : 0;
	3911 : 0;
	3912 : 1;
	3913 : 1;
	3914 : 0;
	3915 : 0;
	3916 : 0;
	3917 : 0;
	3918 : 1;
	3919 : 1;
	3920 : 0;
	3921 : 1;
	3922 : 0;
	3923 : 0;
	3924 : 1;
	3925 : 1;
	3926 : 0;
	3927 : 0;
	3928 : 0;
	3929 : 0;
	3930 : 0;
	3931 : 1;
	3932 : 0;
	3933 : 0;
	3934 : 0;
	3935 : 0;
	3936 : 0;
	3937 : 0;
	3938 : 0;
	3939 : 0;
	3940 : 0;
	3941 : 1;
	3942 : 0;
	3943 : 1;
	3944 : 1;
	3945 : 1;
	3946 : 1;
	3947 : 0;
	3948 : 1;
	3949 : 0;
	3950 : 1;
	3951 : 1;
	3952 : 1;
	3953 : 0;
	3954 : 0;
	3955 : 0;
	3956 : 0;
	3957 : 1;
	3958 : 0;
	3959 : 0;
	3960 : 1;
	3961 : 0;
	3962 : 0;
	3963 : 1;
	3964 : 1;
	3965 : 1;
	3966 : 1;
	3967 : 0;
	3968 : 0;
	3969 : 0;
	3970 : 0;
	3971 : 1;
	3972 : 1;
	3973 : 1;
	3974 : 0;
	3975 : 0;
	3976 : 0;
	3977 : 0;
	3978 : 1;
	3979 : 0;
	3980 : 0;
	3981 : 0;
	3982 : 0;
	3983 : 1;
	3984 : 1;
	3985 : 1;
	3986 : 1;
	3987 : 0;
	3988 : 0;
	3989 : 0;
	3990 : 0;
	3991 : 0;
	3992 : 1;
	3993 : 0;
	3994 : 0;
	3995 : 0;
	3996 : 1;
	3997 : 1;
	3998 : 1;
	3999 : 1;
	4000 : 0;
	4001 : 0;
	4002 : 1;
	4003 : 1;
	4004 : 0;
	4005 : 0;
	4006 : 1;
	4007 : 0;
	4008 : 0;
	4009 : 0;
	4010 : 0;
	4011 : 0;
	4012 : 1;
	4013 : 1;
	4014 : 1;
	4015 : 0;
	4016 : 1;
	4017 : 0;
	4018 : 0;
	4019 : 0;
	4020 : 1;
	4021 : 1;
	4022 : 1;
	4023 : 1;
	4024 : 0;
	4025 : 0;
	4026 : 0;
	4027 : 0;
	4028 : 1;
	4029 : 1;
	4030 : 0;
	4031 : 1;
	4032 : 1;
	4033 : 1;
	4034 : 1;
	4035 : 1;
	4036 : 0;
	4037 : 0;
	4038 : 0;
	4039 : 0;
	4040 : 0;
	4041 : 1;
	4042 : 1;
	4043 : 1;
	4044 : 1;
	4045 : 1;
	4046 : 1;
	4047 : 0;
	4048 : 0;
	4049 : 0;
	4050 : 1;
	4051 : 1;
	4052 : 0;
	4053 : 0;
	4054 : 0;
	4055 : 0;
	4056 : 1;
	4057 : 1;
	4058 : 0;
	4059 : 0;
	4060 : 0;
	4061 : 0;
	4062 : 1;
	4063 : 1;
	4064 : 1;
	4065 : 1;
	4066 : 1;
	4067 : 1;
	4068 : 1;
	4069 : 1;
	4070 : 1;
	4071 : 1;
	4072 : 1;
	4073 : 1;
	4074 : 1;
	4075 : 1;
	4076 : 1;
	4077 : 1;
	4078 : 1;
	4079 : 1;
	4080 : 1;
	4081 : 1;
	4082 : 1;
	4083 : 1;
	4084 : 1;
	4085 : 1;
	4086 : 1;
	4087 : 1;
	4088 : 1;
	4089 : 1;
	4090 : 1;
	4091 : 1;
	4092 : 1;
	4093 : 1;
	4094 : 1;
	4095 : 1;
	4096 : 0;
	4097 : 0;
	4098 : 1;
	4099 : 1;
	4100 : 0;
	4101 : 0;
	4102 : 1;
	4103 : 0;
	4104 : 0;
	4105 : 1;
	4106 : 1;
	4107 : 0;
	4108 : 1;
	4109 : 1;
	4110 : 1;
	4111 : 0;
	4112 : 1;
	4113 : 1;
	4114 : 0;
	4115 : 1;
	4116 : 1;
	4117 : 1;
	4118 : 0;
	4119 : 1;
	4120 : 1;
	4121 : 0;
	4122 : 0;
	4123 : 1;
	4124 : 1;
	4125 : 1;
	4126 : 1;
	4127 : 1;
	4128 : 1;
	4129 : 1;
	4130 : 1;
	4131 : 1;
	4132 : 1;
	4133 : 1;
	4134 : 1;
	4135 : 1;
	4136 : 0;
	4137 : 1;
	4138 : 1;
	4139 : 1;
	4140 : 1;
	4141 : 1;
	4142 : 0;
	4143 : 1;
	4144 : 1;
	4145 : 1;
	4146 : 0;
	4147 : 0;
	4148 : 0;
	4149 : 0;
	4150 : 1;
	4151 : 0;
	4152 : 0;
	4153 : 1;
	4154 : 0;
	4155 : 1;
	4156 : 1;
	4157 : 1;
	4158 : 0;
	4159 : 1;
	4160 : 0;
	4161 : 0;
	4162 : 1;
	4163 : 1;
	4164 : 1;
	4165 : 0;
	4166 : 1;
	4167 : 1;
	4168 : 1;
	4169 : 0;
	4170 : 0;
	4171 : 1;
	4172 : 0;
	4173 : 0;
	4174 : 1;
	4175 : 1;
	4176 : 0;
	4177 : 0;
	4178 : 1;
	4179 : 1;
	4180 : 1;
	4181 : 1;
	4182 : 0;
	4183 : 1;
	4184 : 1;
	4185 : 1;
	4186 : 1;
	4187 : 1;
	4188 : 0;
	4189 : 1;
	4190 : 1;
	4191 : 1;
	4192 : 0;
	4193 : 1;
	4194 : 1;
	4195 : 1;
	4196 : 0;
	4197 : 0;
	4198 : 0;
	4199 : 0;
	4200 : 1;
	4201 : 0;
	4202 : 0;
	4203 : 1;
	4204 : 1;
	4205 : 1;
	4206 : 1;
	4207 : 0;
	4208 : 1;
	4209 : 1;
	4210 : 1;
	4211 : 0;
	4212 : 1;
	4213 : 0;
	4214 : 1;
	4215 : 1;
	4216 : 1;
	4217 : 0;
	4218 : 1;
	4219 : 1;
	4220 : 0;
	4221 : 1;
	4222 : 1;
	4223 : 1;
	4224 : 1;
	4225 : 1;
	4226 : 0;
	4227 : 0;
	4228 : 1;
	4229 : 1;
	4230 : 1;
	4231 : 0;
	4232 : 1;
	4233 : 0;
	4234 : 1;
	4235 : 1;
	4236 : 0;
	4237 : 1;
	4238 : 1;
	4239 : 1;
	4240 : 0;
	4241 : 0;
	4242 : 0;
	4243 : 0;
	4244 : 0;
	4245 : 0;
	4246 : 1;
	4247 : 1;
	4248 : 0;
	4249 : 0;
	4250 : 1;
	4251 : 1;
	4252 : 1;
	4253 : 1;
	4254 : 1;
	4255 : 0;
	4256 : 1;
	4257 : 0;
	4258 : 1;
	4259 : 1;
	4260 : 0;
	4261 : 1;
	4262 : 1;
	4263 : 1;
	4264 : 0;
	4265 : 1;
	4266 : 1;
	4267 : 1;
	4268 : 1;
	4269 : 1;
	4270 : 0;
	4271 : 1;
	4272 : 1;
	4273 : 1;
	4274 : 1;
	4275 : 1;
	4276 : 0;
	4277 : 0;
	4278 : 1;
	4279 : 1;
	4280 : 1;
	4281 : 1;
	4282 : 1;
	4283 : 1;
	4284 : 1;
	4285 : 1;
	4286 : 1;
	4287 : 1;
	4288 : 1;
	4289 : 0;
	4290 : 1;
	4291 : 0;
	4292 : 1;
	4293 : 1;
	4294 : 1;
	4295 : 0;
	4296 : 0;
	4297 : 1;
	4298 : 1;
	4299 : 1;
	4300 : 1;
	4301 : 1;
	4302 : 0;
	4303 : 1;
	4304 : 1;
	4305 : 1;
	4306 : 1;
	4307 : 1;
	4308 : 1;
	4309 : 1;
	4310 : 1;
	4311 : 1;
	4312 : 1;
	4313 : 1;
	4314 : 1;
	4315 : 1;
	4316 : 1;
	4317 : 1;
	4318 : 1;
	4319 : 1;
	4320 : 1;
	4321 : 1;
	4322 : 1;
	4323 : 1;
	4324 : 1;
	4325 : 1;
	4326 : 1;
	4327 : 1;
	4328 : 1;
	4329 : 1;
	4330 : 1;
	4331 : 1;
	4332 : 1;
	4333 : 1;
	4334 : 1;
	4335 : 0;
	4336 : 1;
	4337 : 1;
	4338 : 1;
	4339 : 1;
	4340 : 0;
	4341 : 0;
	4342 : 1;
	4343 : 0;
	4344 : 0;
	4345 : 1;
	4346 : 1;
	4347 : 0;
	4348 : 1;
	4349 : 1;
	4350 : 1;
	4351 : 0;
	4352 : 1;
	4353 : 1;
	4354 : 0;
	4355 : 1;
	4356 : 1;
	4357 : 1;
	4358 : 0;
	4359 : 1;
	4360 : 1;
	4361 : 0;
	4362 : 0;
	4363 : 1;
	4364 : 0;
	4365 : 0;
	4366 : 0;
	4367 : 1;
	4368 : 1;
	4369 : 1;
	4370 : 1;
	4371 : 1;
	4372 : 1;
	4373 : 1;
	4374 : 1;
	4375 : 1;
	4376 : 0;
	4377 : 1;
	4378 : 1;
	4379 : 1;
	4380 : 1;
	4381 : 1;
	4382 : 0;
	4383 : 1;
	4384 : 1;
	4385 : 1;
	4386 : 0;
	4387 : 0;
	4388 : 0;
	4389 : 0;
	4390 : 1;
	4391 : 0;
	4392 : 0;
	4393 : 1;
	4394 : 0;
	4395 : 1;
	4396 : 1;
	4397 : 1;
	4398 : 0;
	4399 : 1;
	4400 : 0;
	4401 : 1;
	4402 : 1;
	4403 : 1;
	4404 : 1;
	4405 : 0;
	4406 : 1;
	4407 : 1;
	4408 : 1;
	4409 : 0;
	4410 : 0;
	4411 : 1;
	4412 : 0;
	4413 : 0;
	4414 : 1;
	4415 : 1;
	4416 : 1;
	4417 : 0;
	4418 : 0;
	4419 : 0;
	4420 : 1;
	4421 : 1;
	4422 : 1;
	4423 : 1;
	4424 : 1;
	4425 : 1;
	4426 : 1;
	4427 : 1;
	4428 : 0;
	4429 : 1;
	4430 : 1;
	4431 : 1;
	4432 : 0;
	4433 : 1;
	4434 : 1;
	4435 : 1;
	4436 : 0;
	4437 : 0;
	4438 : 0;
	4439 : 0;
	4440 : 1;
	4441 : 0;
	4442 : 0;
	4443 : 1;
	4444 : 1;
	4445 : 1;
	4446 : 1;
	4447 : 0;
	4448 : 1;
	4449 : 1;
	4450 : 1;
	4451 : 0;
	4452 : 1;
	4453 : 0;
	4454 : 0;
	4455 : 0;
	4456 : 0;
	4457 : 0;
	4458 : 1;
	4459 : 1;
	4460 : 0;
	4461 : 1;
	4462 : 1;
	4463 : 1;
	4464 : 1;
	4465 : 1;
	4466 : 0;
	4467 : 0;
	4468 : 1;
	4469 : 1;
	4470 : 1;
	4471 : 0;
	4472 : 1;
	4473 : 0;
	4474 : 1;
	4475 : 1;
	4476 : 0;
	4477 : 1;
	4478 : 1;
	4479 : 1;
	4480 : 0;
	4481 : 1;
	4482 : 1;
	4483 : 1;
	4484 : 0;
	4485 : 0;
	4486 : 1;
	4487 : 1;
	4488 : 0;
	4489 : 0;
	4490 : 1;
	4491 : 1;
	4492 : 1;
	4493 : 1;
	4494 : 1;
	4495 : 0;
	4496 : 1;
	4497 : 0;
	4498 : 1;
	4499 : 1;
	4500 : 0;
	4501 : 1;
	4502 : 1;
	4503 : 1;
	4504 : 0;
	4505 : 1;
	4506 : 1;
	4507 : 1;
	4508 : 1;
	4509 : 1;
	4510 : 0;
	4511 : 1;
	4512 : 1;
	4513 : 1;
	4514 : 1;
	4515 : 1;
	4516 : 0;
	4517 : 0;
	4518 : 1;
	4519 : 1;
	4520 : 1;
	4521 : 1;
	4522 : 1;
	4523 : 1;
	4524 : 1;
	4525 : 1;
	4526 : 1;
	4527 : 1;
	4528 : 1;
	4529 : 0;
	4530 : 1;
	4531 : 0;
	4532 : 1;
	4533 : 1;
	4534 : 1;
	4535 : 0;
	4536 : 0;
	4537 : 1;
	4538 : 1;
	4539 : 1;
	4540 : 1;
	4541 : 1;
	4542 : 0;
	4543 : 1;
	4544 : 1;
	4545 : 1;
	4546 : 1;
	4547 : 1;
	4548 : 1;
	4549 : 1;
	4550 : 1;
	4551 : 1;
	4552 : 1;
	4553 : 1;
	4554 : 1;
	4555 : 1;
	4556 : 1;
	4557 : 1;
	4558 : 1;
	4559 : 1;
	4560 : 1;
	4561 : 1;
	4562 : 1;
	4563 : 1;
	4564 : 1;
	4565 : 1;
	4566 : 1;
	4567 : 1;
	4568 : 1;
	4569 : 1;
	4570 : 1;
	4571 : 1;
	4572 : 1;
	4573 : 1;
	4574 : 0;
	4575 : 1;
	4576 : 1;
	4577 : 1;
	4578 : 1;
	4579 : 1;
	4580 : 0;
	4581 : 0;
	4582 : 1;
	4583 : 0;
	4584 : 0;
	4585 : 1;
	4586 : 1;
	4587 : 0;
	4588 : 1;
	4589 : 1;
	4590 : 1;
	4591 : 0;
	4592 : 1;
	4593 : 1;
	4594 : 0;
	4595 : 1;
	4596 : 1;
	4597 : 1;
	4598 : 0;
	4599 : 1;
	4600 : 1;
	4601 : 0;
	4602 : 0;
	4603 : 1;
	4604 : 0;
	4605 : 0;
	4606 : 0;
	4607 : 1;
	4608 : 1;
	4609 : 1;
	4610 : 1;
	4611 : 1;
	4612 : 1;
	4613 : 1;
	4614 : 1;
	4615 : 1;
	4616 : 0;
	4617 : 1;
	4618 : 1;
	4619 : 1;
	4620 : 0;
	4621 : 1;
	4622 : 0;
	4623 : 1;
	4624 : 1;
	4625 : 1;
	4626 : 0;
	4627 : 0;
	4628 : 0;
	4629 : 0;
	4630 : 1;
	4631 : 0;
	4632 : 0;
	4633 : 1;
	4634 : 0;
	4635 : 1;
	4636 : 1;
	4637 : 1;
	4638 : 0;
	4639 : 1;
	4640 : 0;
	4641 : 1;
	4642 : 1;
	4643 : 1;
	4644 : 1;
	4645 : 0;
	4646 : 1;
	4647 : 1;
	4648 : 0;
	4649 : 0;
	4650 : 0;
	4651 : 1;
	4652 : 0;
	4653 : 0;
	4654 : 1;
	4655 : 1;
	4656 : 1;
	4657 : 1;
	4658 : 1;
	4659 : 0;
	4660 : 0;
	4661 : 1;
	4662 : 0;
	4663 : 1;
	4664 : 1;
	4665 : 1;
	4666 : 1;
	4667 : 1;
	4668 : 0;
	4669 : 1;
	4670 : 1;
	4671 : 1;
	4672 : 0;
	4673 : 1;
	4674 : 1;
	4675 : 1;
	4676 : 0;
	4677 : 0;
	4678 : 0;
	4679 : 0;
	4680 : 1;
	4681 : 0;
	4682 : 0;
	4683 : 1;
	4684 : 1;
	4685 : 1;
	4686 : 1;
	4687 : 0;
	4688 : 1;
	4689 : 1;
	4690 : 1;
	4691 : 0;
	4692 : 1;
	4693 : 0;
	4694 : 1;
	4695 : 1;
	4696 : 1;
	4697 : 1;
	4698 : 1;
	4699 : 1;
	4700 : 0;
	4701 : 1;
	4702 : 1;
	4703 : 1;
	4704 : 1;
	4705 : 1;
	4706 : 0;
	4707 : 0;
	4708 : 1;
	4709 : 0;
	4710 : 0;
	4711 : 0;
	4712 : 1;
	4713 : 0;
	4714 : 1;
	4715 : 1;
	4716 : 0;
	4717 : 1;
	4718 : 1;
	4719 : 1;
	4720 : 0;
	4721 : 1;
	4722 : 1;
	4723 : 1;
	4724 : 0;
	4725 : 0;
	4726 : 1;
	4727 : 1;
	4728 : 1;
	4729 : 1;
	4730 : 1;
	4731 : 1;
	4732 : 1;
	4733 : 1;
	4734 : 1;
	4735 : 0;
	4736 : 1;
	4737 : 0;
	4738 : 1;
	4739 : 1;
	4740 : 0;
	4741 : 1;
	4742 : 1;
	4743 : 1;
	4744 : 0;
	4745 : 1;
	4746 : 1;
	4747 : 1;
	4748 : 1;
	4749 : 1;
	4750 : 0;
	4751 : 1;
	4752 : 1;
	4753 : 1;
	4754 : 0;
	4755 : 0;
	4756 : 0;
	4757 : 0;
	4758 : 1;
	4759 : 1;
	4760 : 1;
	4761 : 1;
	4762 : 1;
	4763 : 1;
	4764 : 1;
	4765 : 0;
	4766 : 1;
	4767 : 1;
	4768 : 1;
	4769 : 0;
	4770 : 1;
	4771 : 0;
	4772 : 1;
	4773 : 1;
	4774 : 1;
	4775 : 0;
	4776 : 0;
	4777 : 0;
	4778 : 0;
	4779 : 1;
	4780 : 1;
	4781 : 1;
	4782 : 0;
	4783 : 1;
	4784 : 1;
	4785 : 1;
	4786 : 1;
	4787 : 1;
	4788 : 1;
	4789 : 1;
	4790 : 1;
	4791 : 1;
	4792 : 1;
	4793 : 1;
	4794 : 1;
	4795 : 1;
	4796 : 1;
	4797 : 1;
	4798 : 1;
	4799 : 1;
	4800 : 1;
	4801 : 1;
	4802 : 1;
	4803 : 1;
	4804 : 1;
	4805 : 1;
	4806 : 1;
	4807 : 1;
	4808 : 1;
	4809 : 1;
	4810 : 1;
	4811 : 1;
	4812 : 1;
	4813 : 1;
	4814 : 0;
	4815 : 0;
	4816 : 0;
	4817 : 0;
	4818 : 0;
	4819 : 0;
	4820 : 1;
	4821 : 0;
	4822 : 0;
	4823 : 0;
	4824 : 1;
	4825 : 0;
	4826 : 1;
	4827 : 1;
	4828 : 0;
	4829 : 0;
	4830 : 0;
	4831 : 1;
	4832 : 1;
	4833 : 1;
	4834 : 0;
	4835 : 1;
	4836 : 1;
	4837 : 1;
	4838 : 1;
	4839 : 0;
	4840 : 0;
	4841 : 0;
	4842 : 0;
	4843 : 0;
	4844 : 1;
	4845 : 1;
	4846 : 1;
	4847 : 1;
	4848 : 1;
	4849 : 1;
	4850 : 1;
	4851 : 1;
	4852 : 1;
	4853 : 1;
	4854 : 1;
	4855 : 1;
	4856 : 1;
	4857 : 0;
	4858 : 0;
	4859 : 0;
	4860 : 1;
	4861 : 1;
	4862 : 1;
	4863 : 0;
	4864 : 0;
	4865 : 0;
	4866 : 0;
	4867 : 1;
	4868 : 0;
	4869 : 0;
	4870 : 1;
	4871 : 0;
	4872 : 0;
	4873 : 1;
	4874 : 1;
	4875 : 0;
	4876 : 0;
	4877 : 0;
	4878 : 0;
	4879 : 1;
	4880 : 0;
	4881 : 1;
	4882 : 1;
	4883 : 1;
	4884 : 1;
	4885 : 1;
	4886 : 0;
	4887 : 0;
	4888 : 0;
	4889 : 0;
	4890 : 0;
	4891 : 1;
	4892 : 0;
	4893 : 0;
	4894 : 0;
	4895 : 0;
	4896 : 0;
	4897 : 0;
	4898 : 0;
	4899 : 0;
	4900 : 0;
	4901 : 1;
	4902 : 0;
	4903 : 1;
	4904 : 1;
	4905 : 1;
	4906 : 1;
	4907 : 1;
	4908 : 0;
	4909 : 1;
	4910 : 1;
	4911 : 1;
	4912 : 1;
	4913 : 0;
	4914 : 0;
	4915 : 0;
	4916 : 0;
	4917 : 1;
	4918 : 1;
	4919 : 0;
	4920 : 0;
	4921 : 0;
	4922 : 1;
	4923 : 0;
	4924 : 1;
	4925 : 1;
	4926 : 1;
	4927 : 1;
	4928 : 0;
	4929 : 0;
	4930 : 0;
	4931 : 0;
	4932 : 1;
	4933 : 1;
	4934 : 0;
	4935 : 0;
	4936 : 0;
	4937 : 0;
	4938 : 1;
	4939 : 1;
	4940 : 0;
	4941 : 0;
	4942 : 0;
	4943 : 0;
	4944 : 1;
	4945 : 1;
	4946 : 1;
	4947 : 0;
	4948 : 0;
	4949 : 0;
	4950 : 1;
	4951 : 0;
	4952 : 1;
	4953 : 0;
	4954 : 1;
	4955 : 1;
	4956 : 0;
	4957 : 1;
	4958 : 1;
	4959 : 1;
	4960 : 0;
	4961 : 1;
	4962 : 1;
	4963 : 1;
	4964 : 0;
	4965 : 0;
	4966 : 1;
	4967 : 1;
	4968 : 1;
	4969 : 1;
	4970 : 1;
	4971 : 1;
	4972 : 1;
	4973 : 1;
	4974 : 1;
	4975 : 0;
	4976 : 1;
	4977 : 0;
	4978 : 1;
	4979 : 1;
	4980 : 0;
	4981 : 1;
	4982 : 1;
	4983 : 1;
	4984 : 0;
	4985 : 0;
	4986 : 0;
	4987 : 0;
	4988 : 0;
	4989 : 1;
	4990 : 1;
	4991 : 0;
	4992 : 0;
	4993 : 0;
	4994 : 0;
	4995 : 1;
	4996 : 0;
	4997 : 0;
	4998 : 0;
	4999 : 0;
	5000 : 0;
	5001 : 0;
	5002 : 1;
	5003 : 1;
	5004 : 1;
	5005 : 1;
	5006 : 0;
	5007 : 0;
	5008 : 0;
	5009 : 1;
	5010 : 1;
	5011 : 1;
	5012 : 0;
	5013 : 0;
	5014 : 0;
	5015 : 0;
	5016 : 1;
	5017 : 1;
	5018 : 0;
	5019 : 0;
	5020 : 0;
	5021 : 0;
	5022 : 1;
	5023 : 1;
	5024 : 1;
	5025 : 1;
	5026 : 1;
	5027 : 1;
	5028 : 1;
	5029 : 1;
	5030 : 1;
	5031 : 1;
	5032 : 1;
	5033 : 1;
	5034 : 1;
	5035 : 1;
	5036 : 1;
	5037 : 1;
	5038 : 1;
	5039 : 1;
	5040 : 1;
	5041 : 1;
	5042 : 1;
	5043 : 1;
	5044 : 1;
	5045 : 1;
	5046 : 1;
	5047 : 1;
	5048 : 1;
	5049 : 1;
	5050 : 1;
	5051 : 1;
	5052 : 1;
	5053 : 1;
	5054 : 1;
	5055 : 1;
	5056 : 1;
	5057 : 1;
	5058 : 1;
	5059 : 1;
	5060 : 1;
	5061 : 1;
	5062 : 1;
	5063 : 1;
	5064 : 1;
	5065 : 1;
	5066 : 1;
	5067 : 1;
	5068 : 1;
	5069 : 1;
	5070 : 1;
	5071 : 1;
	5072 : 1;
	5073 : 1;
	5074 : 1;
	5075 : 1;
	5076 : 1;
	5077 : 1;
	5078 : 1;
	5079 : 1;
	5080 : 1;
	5081 : 1;
	5082 : 1;
	5083 : 1;
	5084 : 1;
	5085 : 1;
	5086 : 1;
	5087 : 1;
	5088 : 1;
	5089 : 1;
	5090 : 1;
	5091 : 1;
	5092 : 1;
	5093 : 1;
	5094 : 1;
	5095 : 1;
	5096 : 1;
	5097 : 1;
	5098 : 1;
	5099 : 1;
	5100 : 1;
	5101 : 1;
	5102 : 1;
	5103 : 1;
	5104 : 1;
	5105 : 1;
	5106 : 1;
	5107 : 1;
	5108 : 1;
	5109 : 1;
	5110 : 1;
	5111 : 1;
	5112 : 1;
	5113 : 1;
	5114 : 1;
	5115 : 1;
	5116 : 1;
	5117 : 1;
	5118 : 0;
	5119 : 1;
	5120 : 1;
	5121 : 1;
	5122 : 1;
	5123 : 1;
	5124 : 1;
	5125 : 1;
	5126 : 1;
	5127 : 1;
	5128 : 1;
	5129 : 1;
	5130 : 1;
	5131 : 1;
	5132 : 1;
	5133 : 1;
	5134 : 1;
	5135 : 1;
	5136 : 1;
	5137 : 1;
	5138 : 1;
	5139 : 1;
	5140 : 1;
	5141 : 1;
	5142 : 1;
	5143 : 1;
	5144 : 1;
	5145 : 1;
	5146 : 1;
	5147 : 1;
	5148 : 1;
	5149 : 1;
	5150 : 1;
	5151 : 1;
	5152 : 1;
	5153 : 1;
	5154 : 1;
	5155 : 1;
	5156 : 1;
	5157 : 1;
	5158 : 1;
	5159 : 1;
	5160 : 1;
	5161 : 1;
	5162 : 1;
	5163 : 1;
	5164 : 1;
	5165 : 1;
	5166 : 1;
	5167 : 1;
	5168 : 1;
	5169 : 1;
	5170 : 1;
	5171 : 0;
	5172 : 1;
	5173 : 1;
	5174 : 1;
	5175 : 1;
	5176 : 1;
	5177 : 1;
	5178 : 1;
	5179 : 1;
	5180 : 1;
	5181 : 1;
	5182 : 1;
	5183 : 1;
	5184 : 1;
	5185 : 1;
	5186 : 1;
	5187 : 1;
	5188 : 1;
	5189 : 1;
	5190 : 1;
	5191 : 1;
	5192 : 1;
	5193 : 1;
	5194 : 1;
	5195 : 1;
	5196 : 1;
	5197 : 1;
	5198 : 1;
	5199 : 1;
	5200 : 1;
	5201 : 1;
	5202 : 1;
	5203 : 1;
	5204 : 1;
	5205 : 1;
	5206 : 1;
	5207 : 1;
	5208 : 1;
	5209 : 1;
	5210 : 1;
	5211 : 1;
	5212 : 1;
	5213 : 1;
	5214 : 1;
	5215 : 1;
	5216 : 1;
	5217 : 1;
	5218 : 1;
	5219 : 1;
	5220 : 1;
	5221 : 1;
	5222 : 1;
	5223 : 1;
	5224 : 1;
	5225 : 1;
	5226 : 1;
	5227 : 1;
	5228 : 1;
	5229 : 1;
	5230 : 1;
	5231 : 1;
	5232 : 1;
	5233 : 1;
	5234 : 1;
	5235 : 1;
	5236 : 1;
	5237 : 1;
	5238 : 1;
	5239 : 1;
	5240 : 1;
	5241 : 1;
	5242 : 1;
	5243 : 1;
	5244 : 1;
	5245 : 1;
	5246 : 1;
	5247 : 1;
	5248 : 1;
	5249 : 1;
	5250 : 1;
	5251 : 1;
	5252 : 1;
	5253 : 1;
	5254 : 1;
	5255 : 1;
	5256 : 1;
	5257 : 1;
	5258 : 1;
	5259 : 1;
	5260 : 1;
	5261 : 1;
	5262 : 1;
	5263 : 1;
	5264 : 1;
	5265 : 1;
	5266 : 1;
	5267 : 1;
	5268 : 1;
	5269 : 1;
	5270 : 1;
	5271 : 1;
	5272 : 1;
	5273 : 1;
	5274 : 1;
	5275 : 1;
	5276 : 1;
	5277 : 1;
	5278 : 1;
	5279 : 1;
	5280 : 1;
	5281 : 1;
	5282 : 1;
	5283 : 1;
	5284 : 1;
	5285 : 1;
	5286 : 1;
	5287 : 1;
	5288 : 1;
	5289 : 1;
	5290 : 1;
	5291 : 1;
	5292 : 1;
	5293 : 1;
	5294 : 1;
	5295 : 1;
	5296 : 1;
	5297 : 1;
	5298 : 1;
	5299 : 1;
	5300 : 1;
	5301 : 1;
	5302 : 1;
	5303 : 1;
	5304 : 1;
	5305 : 1;
	5306 : 1;
	5307 : 1;
	5308 : 1;
	5309 : 1;
	5310 : 1;
	5311 : 1;
	5312 : 1;
	5313 : 1;
	5314 : 1;
	5315 : 1;
	5316 : 1;
	5317 : 1;
	5318 : 1;
	5319 : 1;
	5320 : 1;
	5321 : 1;
	5322 : 1;
	5323 : 1;
	5324 : 1;
	5325 : 1;
	5326 : 1;
	5327 : 1;
	5328 : 1;
	5329 : 1;
	5330 : 1;
	5331 : 1;
	5332 : 1;
	5333 : 1;
	5334 : 1;
	5335 : 1;
	5336 : 1;
	5337 : 1;
	5338 : 1;
	5339 : 1;
	5340 : 1;
	5341 : 1;
	5342 : 1;
	5343 : 1;
	5344 : 1;
	5345 : 1;
	5346 : 1;
	5347 : 1;
	5348 : 1;
	5349 : 1;
	5350 : 1;
	5351 : 1;
	5352 : 1;
	5353 : 1;
	5354 : 1;
	5355 : 0;
	5356 : 0;
	5357 : 0;
	5358 : 1;
	5359 : 1;
	5360 : 1;
	5361 : 1;
	5362 : 1;
	5363 : 1;
	5364 : 1;
	5365 : 1;
	5366 : 1;
	5367 : 1;
	5368 : 1;
	5369 : 1;
	5370 : 1;
	5371 : 1;
	5372 : 1;
	5373 : 1;
	5374 : 1;
	5375 : 1;
	5376 : 1;
	5377 : 1;
	5378 : 1;
	5379 : 1;
	5380 : 1;
	5381 : 1;
	5382 : 1;
	5383 : 1;
	5384 : 1;
	5385 : 1;
	5386 : 1;
	5387 : 1;
	5388 : 1;
	5389 : 1;
	5390 : 1;
	5391 : 1;
	5392 : 1;
	5393 : 1;
	5394 : 1;
	5395 : 1;
	5396 : 1;
	5397 : 1;
	5398 : 1;
	5399 : 1;
	5400 : 1;
	5401 : 1;
	5402 : 1;
	5403 : 1;
	5404 : 1;
	5405 : 1;
	5406 : 1;
	5407 : 1;
	5408 : 0;
	5409 : 0;
	5410 : 0;
	5411 : 1;
	5412 : 1;
	5413 : 1;
	5414 : 1;
	5415 : 1;
	5416 : 1;
	5417 : 1;
	5418 : 1;
	5419 : 1;
	5420 : 1;
	5421 : 1;
	5422 : 1;
	5423 : 1;
	5424 : 1;
	5425 : 1;
	5426 : 1;
	5427 : 1;
	5428 : 1;
	5429 : 1;
	5430 : 1;
	5431 : 1;
	5432 : 1;
	5433 : 1;
	5434 : 1;
	5435 : 1;
	5436 : 1;
	5437 : 1;
	5438 : 1;
	5439 : 1;
	5440 : 1;
	5441 : 1;
	5442 : 1;
	5443 : 1;
	5444 : 1;
	5445 : 1;
	5446 : 1;
	5447 : 1;
	5448 : 1;
	5449 : 1;
	5450 : 1;
	5451 : 1;
	5452 : 1;
	5453 : 1;
	5454 : 1;
	5455 : 1;
	5456 : 1;
	5457 : 1;
	5458 : 1;
	5459 : 1;
	5460 : 1;
	5461 : 1;
	5462 : 1;
	5463 : 1;
	5464 : 1;
	5465 : 1;
	5466 : 1;
	5467 : 1;
	5468 : 1;
	5469 : 1;
	5470 : 1;
	5471 : 1;
	5472 : 1;
	5473 : 1;
	5474 : 1;
	5475 : 1;
	5476 : 1;
	5477 : 1;
	5478 : 1;
	5479 : 1;
	5480 : 1;
	5481 : 1;
	5482 : 1;
	5483 : 1;
	5484 : 1;
	5485 : 1;
	5486 : 1;
	5487 : 1;
	5488 : 1;
	5489 : 1;
	5490 : 1;
	5491 : 1;
	5492 : 1;
	5493 : 1;
	5494 : 1;
	5495 : 1;
	5496 : 1;
	5497 : 1;
	5498 : 1;
	5499 : 1;
	5500 : 1;
	5501 : 1;
	5502 : 1;
	5503 : 1;
	5504 : 1;
	5505 : 1;
	5506 : 1;
	5507 : 1;
	5508 : 1;
	5509 : 1;
	5510 : 1;
	5511 : 1;
	5512 : 1;
	5513 : 1;
	5514 : 1;
	5515 : 1;
	5516 : 1;
	5517 : 1;
	5518 : 1;
	5519 : 1;
	5520 : 1;
	5521 : 1;
	5522 : 1;
	5523 : 1;
	5524 : 1;
	5525 : 1;
	5526 : 1;
	5527 : 1;
	5528 : 1;
	5529 : 1;
	5530 : 1;
	5531 : 1;
	5532 : 1;
	5533 : 1;
	5534 : 1;
	5535 : 1;
	5536 : 1;
	5537 : 1;
	5538 : 1;
	5539 : 1;
	5540 : 1;
	5541 : 1;
	5542 : 1;
	5543 : 1;
	5544 : 1;
	5545 : 1;
	5546 : 1;
	5547 : 1;
	5548 : 1;
	5549 : 1;
	5550 : 1;
	5551 : 1;
	5552 : 1;
	5553 : 1;
	5554 : 1;
	5555 : 1;
	5556 : 1;
	5557 : 1;
	5558 : 1;
	5559 : 1;
	5560 : 1;
	5561 : 1;
	5562 : 1;
	5563 : 1;
	5564 : 1;
	5565 : 1;
	5566 : 1;
	5567 : 1;
	5568 : 1;
	5569 : 1;
	5570 : 1;
	5571 : 1;
	5572 : 1;
	5573 : 1;
	5574 : 1;
	5575 : 1;
	5576 : 1;
	5577 : 1;
	5578 : 1;
	5579 : 1;
	5580 : 1;
	5581 : 1;
	5582 : 1;
	5583 : 1;
	5584 : 1;
	5585 : 1;
	5586 : 1;
	5587 : 1;
	5588 : 1;
	5589 : 1;
	5590 : 1;
	5591 : 1;
	5592 : 1;
	5593 : 1;
	5594 : 1;
	5595 : 1;
	5596 : 1;
	5597 : 1;
	5598 : 1;
	5599 : 1;
	5600 : 1;
	5601 : 1;
	5602 : 1;
	5603 : 1;
	5604 : 1;
	5605 : 1;
	5606 : 1;
	5607 : 1;
	5608 : 1;
	5609 : 1;
	5610 : 1;
	5611 : 1;
	5612 : 1;
	5613 : 1;
	5614 : 1;
	5615 : 1;
	5616 : 1;
	5617 : 1;
	5618 : 1;
	5619 : 1;
	5620 : 1;
	5621 : 1;
	5622 : 1;
	5623 : 1;
	5624 : 1;
	5625 : 1;
	5626 : 1;
	5627 : 1;
	5628 : 1;
	5629 : 1;
	5630 : 1;
	5631 : 1;
	5632 : 1;
	5633 : 1;
	5634 : 1;
	5635 : 1;
	5636 : 1;
	5637 : 1;
	5638 : 1;
	5639 : 1;
	5640 : 1;
	5641 : 1;
	5642 : 1;
	5643 : 1;
	5644 : 1;
	5645 : 1;
	5646 : 1;
	5647 : 1;
	5648 : 1;
	5649 : 1;
	5650 : 1;
	5651 : 1;
	5652 : 1;
	5653 : 1;
	5654 : 1;
	5655 : 1;
	5656 : 1;
	5657 : 1;
	5658 : 1;
	5659 : 1;
	5660 : 1;
	5661 : 1;
	5662 : 1;
	5663 : 1;
	5664 : 1;
	5665 : 1;
	5666 : 1;
	5667 : 1;
	5668 : 1;
	5669 : 1;
	5670 : 1;
	5671 : 1;
	5672 : 1;
	5673 : 1;
	5674 : 1;
	5675 : 1;
	5676 : 1;
	5677 : 1;
	5678 : 1;
	5679 : 1;
	5680 : 1;
	5681 : 1;
	5682 : 1;
	5683 : 1;
	5684 : 1;
	5685 : 1;
	5686 : 1;
	5687 : 1;
	5688 : 1;
	5689 : 1;
	5690 : 1;
	5691 : 1;
	5692 : 1;
	5693 : 1;
	5694 : 1;
	5695 : 1;
	5696 : 1;
	5697 : 1;
	5698 : 1;
	5699 : 1;
	5700 : 1;
	5701 : 1;
	5702 : 1;
	5703 : 1;
	5704 : 1;
	5705 : 1;
	5706 : 1;
	5707 : 1;
	5708 : 1;
	5709 : 1;
	5710 : 1;
	5711 : 1;
	5712 : 1;
	5713 : 1;
	5714 : 1;
	5715 : 1;
	5716 : 1;
	5717 : 1;
	5718 : 1;
	5719 : 1;
	5720 : 1;
	5721 : 1;
	5722 : 1;
	5723 : 1;
	5724 : 1;
	5725 : 1;
	5726 : 1;
	5727 : 1;
	5728 : 1;
	5729 : 1;
	5730 : 1;
	5731 : 1;
	5732 : 1;
	5733 : 1;
	5734 : 1;
	5735 : 1;
	5736 : 1;
	5737 : 1;
	5738 : 1;
	5739 : 1;
	5740 : 1;
	5741 : 1;
	5742 : 1;
	5743 : 1;
	5744 : 1;
	5745 : 1;
	5746 : 1;
	5747 : 1;
	5748 : 1;
	5749 : 1;
	5750 : 1;
	5751 : 1;
	5752 : 1;
	5753 : 1;
	5754 : 1;
	5755 : 1;
	5756 : 1;
	5757 : 1;
	5758 : 1;
	5759 : 1;
	5760 : 1;
	5761 : 1;
	5762 : 1;
	5763 : 1;
	5764 : 1;
	5765 : 1;
	5766 : 1;
	5767 : 1;
	5768 : 1;
	5769 : 1;
	5770 : 1;
	5771 : 1;
	5772 : 1;
	5773 : 1;
	5774 : 1;
	5775 : 1;
	5776 : 1;
	5777 : 1;
	5778 : 1;
	5779 : 1;
	5780 : 1;
	5781 : 1;
	5782 : 1;
	5783 : 1;
	5784 : 1;
	5785 : 1;
	5786 : 1;
	5787 : 1;
	5788 : 1;
	5789 : 1;
	5790 : 1;
	5791 : 1;
	5792 : 1;
	5793 : 1;
	5794 : 1;
	5795 : 1;
	5796 : 1;
	5797 : 1;
	5798 : 1;
	5799 : 1;
	5800 : 1;
	5801 : 1;
	5802 : 1;
	5803 : 1;
	5804 : 1;
	5805 : 1;
	5806 : 1;
	5807 : 1;
	5808 : 1;
	5809 : 1;
	5810 : 1;
	5811 : 1;
	5812 : 1;
	5813 : 1;
	5814 : 1;
	5815 : 1;
	5816 : 1;
	5817 : 1;
	5818 : 1;
	5819 : 1;
	5820 : 1;
	5821 : 1;
	5822 : 1;
	5823 : 1;
	5824 : 1;
	5825 : 1;
	5826 : 1;
	5827 : 1;
	5828 : 1;
	5829 : 1;
	5830 : 1;
	5831 : 1;
	5832 : 1;
	5833 : 1;
	5834 : 1;
	5835 : 1;
	5836 : 1;
	5837 : 1;
	5838 : 1;
	5839 : 1;
	5840 : 1;
	5841 : 1;
	5842 : 1;
	5843 : 1;
	5844 : 1;
	5845 : 1;
	5846 : 1;
	5847 : 1;
	5848 : 1;
	5849 : 1;
	5850 : 1;
	5851 : 1;
	5852 : 1;
	5853 : 1;
	5854 : 1;
	5855 : 1;
	5856 : 1;
	5857 : 1;
	5858 : 1;
	5859 : 1;
	5860 : 1;
	5861 : 1;
	5862 : 1;
	5863 : 1;
	5864 : 1;
	5865 : 1;
	5866 : 1;
	5867 : 1;
	5868 : 1;
	5869 : 1;
	5870 : 1;
	5871 : 1;
	5872 : 1;
	5873 : 1;
	5874 : 1;
	5875 : 1;
	5876 : 1;
	5877 : 1;
	5878 : 1;
	5879 : 1;
	5880 : 1;
	5881 : 1;
	5882 : 1;
	5883 : 1;
	5884 : 1;
	5885 : 1;
	5886 : 1;
	5887 : 1;
	5888 : 1;
	5889 : 1;
	5890 : 1;
	5891 : 1;
	5892 : 1;
	5893 : 1;
	5894 : 1;
	5895 : 1;
	5896 : 1;
	5897 : 1;
	5898 : 1;
	5899 : 1;
	5900 : 1;
	5901 : 1;
	5902 : 1;
	5903 : 1;
	5904 : 1;
	5905 : 1;
	5906 : 1;
	5907 : 1;
	5908 : 1;
	5909 : 1;
	5910 : 1;
	5911 : 1;
	5912 : 1;
	5913 : 1;
	5914 : 1;
	5915 : 1;
	5916 : 1;
	5917 : 1;
	5918 : 1;
	5919 : 1;
	5920 : 1;
	5921 : 1;
	5922 : 1;
	5923 : 1;
	5924 : 1;
	5925 : 1;
	5926 : 1;
	5927 : 1;
	5928 : 1;
	5929 : 1;
	5930 : 1;
	5931 : 1;
	5932 : 1;
	5933 : 1;
	5934 : 1;
	5935 : 1;
	5936 : 1;
	5937 : 1;
	5938 : 1;
	5939 : 1;
	5940 : 1;
	5941 : 1;
	5942 : 1;
	5943 : 1;
	5944 : 1;
	5945 : 1;
	5946 : 1;
	5947 : 1;
	5948 : 1;
	5949 : 1;
	5950 : 1;
	5951 : 1;
	5952 : 1;
	5953 : 1;
	5954 : 1;
	5955 : 1;
	5956 : 1;
	5957 : 1;
	5958 : 1;
	5959 : 1;
	5960 : 1;
	5961 : 1;
	5962 : 1;
	5963 : 1;
	5964 : 1;
	5965 : 1;
	5966 : 1;
	5967 : 1;
	5968 : 1;
	5969 : 1;
	5970 : 1;
	5971 : 1;
	5972 : 1;
	5973 : 1;
	5974 : 1;
	5975 : 1;
	5976 : 1;
	5977 : 1;
	5978 : 1;
	5979 : 1;
	5980 : 1;
	5981 : 1;
	5982 : 1;
	5983 : 1;
	5984 : 1;
	5985 : 1;
	5986 : 1;
	5987 : 1;
	5988 : 1;
	5989 : 1;
	5990 : 1;
	5991 : 1;
	5992 : 1;
	5993 : 1;
	5994 : 1;
	5995 : 1;
	5996 : 1;
	5997 : 1;
	5998 : 1;
	5999 : 1;
	6000 : 1;
	6001 : 1;
	6002 : 1;
	6003 : 1;
	6004 : 1;
	6005 : 1;
	6006 : 1;
	6007 : 1;
	6008 : 1;
	6009 : 1;
	6010 : 1;
	6011 : 1;
	6012 : 1;
	6013 : 1;
	6014 : 1;
	6015 : 1;
	6016 : 1;
	6017 : 1;
	6018 : 1;
	6019 : 1;
	6020 : 1;
	6021 : 1;
	6022 : 1;
	6023 : 1;
	6024 : 1;
	6025 : 1;
	6026 : 1;
	6027 : 1;
	6028 : 1;
	6029 : 1;
	6030 : 1;
	6031 : 1;
	6032 : 1;
	6033 : 1;
	6034 : 1;
	6035 : 1;
	6036 : 1;
	6037 : 1;
	6038 : 1;
	6039 : 1;
	6040 : 1;
	6041 : 1;
	6042 : 1;
	6043 : 1;
	6044 : 1;
	6045 : 1;
	6046 : 1;
	6047 : 1;
	6048 : 1;
	6049 : 1;
	6050 : 1;
	6051 : 1;
	6052 : 1;
	6053 : 1;
	6054 : 1;
	6055 : 1;
	6056 : 1;
	6057 : 1;
	6058 : 1;
	6059 : 1;
	6060 : 1;
	6061 : 1;
	6062 : 1;
	6063 : 1;
	6064 : 1;
	6065 : 1;
	6066 : 1;
	6067 : 1;
	6068 : 1;
	6069 : 1;
	6070 : 1;
	6071 : 1;
	6072 : 1;
	6073 : 1;
	6074 : 1;
	6075 : 1;
	6076 : 1;
	6077 : 1;
	6078 : 1;
	6079 : 1;
	6080 : 1;
	6081 : 1;
	6082 : 1;
	6083 : 1;
	6084 : 1;
	6085 : 1;
	6086 : 1;
	6087 : 1;
	6088 : 1;
	6089 : 1;
	6090 : 1;
	6091 : 1;
	6092 : 1;
	6093 : 1;
	6094 : 1;
	6095 : 1;
	6096 : 1;
	6097 : 1;
	6098 : 1;
	6099 : 1;
	6100 : 1;
	6101 : 1;
	6102 : 1;
	6103 : 1;
	6104 : 1;
	6105 : 1;
	6106 : 1;
	6107 : 1;
	6108 : 1;
	6109 : 1;
	6110 : 1;
	6111 : 1;
	6112 : 1;
	6113 : 1;
	6114 : 1;
	6115 : 1;
	6116 : 1;
	6117 : 1;
	6118 : 1;
	6119 : 1;
	6120 : 1;
	6121 : 1;
	6122 : 1;
	6123 : 1;
	6124 : 1;
	6125 : 1;
	6126 : 1;
	6127 : 1;
	6128 : 1;
	6129 : 1;
	6130 : 1;
	6131 : 1;
	6132 : 1;
	6133 : 1;
	6134 : 1;
	6135 : 1;
	6136 : 1;
	6137 : 1;
	6138 : 1;
	6139 : 1;
	6140 : 1;
	6141 : 1;
	6142 : 1;
	6143 : 1;
	6144 : 1;
	6145 : 1;
	6146 : 1;
	6147 : 1;
	6148 : 1;
	6149 : 1;
	6150 : 1;
	6151 : 1;
	6152 : 1;
	6153 : 1;
	6154 : 1;
	6155 : 1;
	6156 : 1;
	6157 : 1;
	6158 : 1;
	6159 : 1;
	6160 : 1;
	6161 : 1;
	6162 : 1;
	6163 : 1;
	6164 : 1;
	6165 : 1;
	6166 : 1;
	6167 : 1;
	6168 : 1;
	6169 : 1;
	6170 : 1;
	6171 : 1;
	6172 : 1;
	6173 : 1;
	6174 : 1;
	6175 : 1;
	6176 : 1;
	6177 : 1;
	6178 : 1;
	6179 : 1;
	6180 : 1;
	6181 : 1;
	6182 : 1;
	6183 : 1;
	6184 : 1;
	6185 : 1;
	6186 : 1;
	6187 : 1;
	6188 : 1;
	6189 : 1;
	6190 : 1;
	6191 : 1;
	6192 : 1;
	6193 : 1;
	6194 : 1;
	6195 : 1;
	6196 : 1;
	6197 : 1;
	6198 : 1;
	6199 : 1;
	6200 : 1;
	6201 : 1;
	6202 : 1;
	6203 : 1;
	6204 : 1;
	6205 : 1;
	6206 : 1;
	6207 : 1;
	6208 : 1;
	6209 : 1;
	6210 : 1;
	6211 : 1;
	6212 : 1;
	6213 : 1;
	6214 : 1;
	6215 : 1;
	6216 : 1;
	6217 : 1;
	6218 : 1;
	6219 : 1;
	6220 : 1;
	6221 : 1;
	6222 : 1;
	6223 : 1;
	6224 : 1;
	6225 : 1;
	6226 : 1;
	6227 : 1;
	6228 : 1;
	6229 : 1;
	6230 : 1;
	6231 : 1;
	6232 : 1;
	6233 : 1;
	6234 : 1;
	6235 : 1;
	6236 : 1;
	6237 : 1;
	6238 : 1;
	6239 : 1;
	6240 : 1;
	6241 : 1;
	6242 : 1;
	6243 : 1;
	6244 : 1;
	6245 : 1;
	6246 : 1;
	6247 : 1;
	6248 : 1;
	6249 : 1;
	6250 : 1;
	6251 : 1;
	6252 : 1;
	6253 : 1;
	6254 : 1;
	6255 : 1;
	6256 : 1;
	6257 : 1;
	6258 : 1;
	6259 : 1;
	6260 : 1;
	6261 : 1;
	6262 : 1;
	6263 : 1;
	6264 : 1;
	6265 : 1;
	6266 : 1;
	6267 : 1;
	6268 : 1;
	6269 : 1;
	6270 : 1;
	6271 : 1;
	6272 : 1;
	6273 : 1;
	6274 : 1;
	6275 : 1;
	6276 : 1;
	6277 : 1;
	6278 : 1;
	6279 : 1;
	6280 : 1;
	6281 : 1;
	6282 : 1;
	6283 : 1;
	6284 : 1;
	6285 : 1;
	6286 : 1;
	6287 : 1;
	6288 : 1;
	6289 : 1;
	6290 : 1;
	6291 : 1;
	6292 : 1;
	6293 : 1;
	6294 : 1;
	6295 : 1;
	6296 : 1;
	6297 : 1;
	6298 : 1;
	6299 : 1;
	6300 : 1;
	6301 : 1;
	6302 : 1;
	6303 : 1;
	6304 : 1;
	6305 : 1;
	6306 : 1;
	6307 : 1;
	6308 : 1;
	6309 : 1;
	6310 : 1;
	6311 : 1;
	6312 : 1;
	6313 : 1;
	6314 : 1;
	6315 : 1;
	6316 : 1;
	6317 : 1;
	6318 : 1;
	6319 : 1;
	6320 : 1;
	6321 : 1;
	6322 : 1;
	6323 : 1;
	6324 : 1;
	6325 : 1;
	6326 : 1;
	6327 : 1;
	6328 : 1;
	6329 : 1;
	6330 : 1;
	6331 : 1;
	6332 : 1;
	6333 : 1;
	6334 : 1;
	6335 : 1;
	6336 : 1;
	6337 : 1;
	6338 : 1;
	6339 : 1;
	6340 : 1;
	6341 : 1;
	6342 : 1;
	6343 : 1;
	6344 : 1;
	6345 : 1;
	6346 : 1;
	6347 : 1;
	6348 : 1;
	6349 : 1;
	6350 : 1;
	6351 : 1;
	6352 : 1;
	6353 : 1;
	6354 : 1;
	6355 : 1;
	6356 : 1;
	6357 : 1;
	6358 : 1;
	6359 : 1;
	6360 : 1;
	6361 : 1;
	6362 : 1;
	6363 : 1;
	6364 : 1;
	6365 : 1;
	6366 : 1;
	6367 : 1;
	6368 : 1;
	6369 : 1;
	6370 : 1;
	6371 : 1;
	6372 : 1;
	6373 : 1;
	6374 : 1;
	6375 : 1;
	6376 : 1;
	6377 : 1;
	6378 : 1;
	6379 : 1;
	6380 : 1;
	6381 : 1;
	6382 : 1;
	6383 : 1;
	6384 : 1;
	6385 : 1;
	6386 : 1;
	6387 : 1;
	6388 : 1;
	6389 : 1;
	6390 : 1;
	6391 : 1;
	6392 : 1;
	6393 : 1;
	6394 : 1;
	6395 : 1;
	6396 : 1;
	6397 : 1;
	6398 : 1;
	6399 : 1;
	6400 : 1;
	6401 : 1;
	6402 : 1;
	6403 : 1;
	6404 : 1;
	6405 : 1;
	6406 : 1;
	6407 : 1;
	6408 : 1;
	6409 : 1;
	6410 : 1;
	6411 : 1;
	6412 : 1;
	6413 : 1;
	6414 : 1;
	6415 : 1;
	6416 : 1;
	6417 : 1;
	6418 : 1;
	6419 : 1;
	6420 : 1;
	6421 : 1;
	6422 : 1;
	6423 : 1;
	6424 : 1;
	6425 : 1;
	6426 : 1;
	6427 : 1;
	6428 : 1;
	6429 : 1;
	6430 : 1;
	6431 : 1;
	6432 : 1;
	6433 : 1;
	6434 : 1;
	6435 : 1;
	6436 : 1;
	6437 : 1;
	6438 : 1;
	6439 : 1;
	6440 : 1;
	6441 : 1;
	6442 : 1;
	6443 : 1;
	6444 : 1;
	6445 : 1;
	6446 : 1;
	6447 : 1;
	6448 : 1;
	6449 : 1;
	6450 : 1;
	6451 : 1;
	6452 : 1;
	6453 : 1;
	6454 : 1;
	6455 : 1;
	6456 : 1;
	6457 : 1;
	6458 : 1;
	6459 : 1;
	6460 : 1;
	6461 : 1;
	6462 : 1;
	6463 : 1;
	6464 : 1;
	6465 : 1;
	6466 : 1;
	6467 : 1;
	6468 : 1;
	6469 : 1;
	6470 : 1;
	6471 : 1;
	6472 : 1;
	6473 : 1;
	6474 : 1;
	6475 : 1;
	6476 : 1;
	6477 : 1;
	6478 : 1;
	6479 : 1;
	6480 : 1;
	6481 : 1;
	6482 : 1;
	6483 : 1;
	6484 : 1;
	6485 : 1;
	6486 : 1;
	6487 : 1;
	6488 : 1;
	6489 : 1;
	6490 : 1;
	6491 : 1;
	6492 : 1;
	6493 : 1;
	6494 : 1;
	6495 : 1;
	6496 : 1;
	6497 : 1;
	6498 : 1;
	6499 : 1;
	6500 : 1;
	6501 : 1;
	6502 : 1;
	6503 : 1;
	6504 : 1;
	6505 : 1;
	6506 : 1;
	6507 : 1;
	6508 : 1;
	6509 : 1;
	6510 : 1;
	6511 : 1;
	6512 : 1;
	6513 : 1;
	6514 : 1;
	6515 : 1;
	6516 : 1;
	6517 : 1;
	6518 : 1;
	6519 : 1;
	6520 : 1;
	6521 : 1;
	6522 : 1;
	6523 : 1;
	6524 : 1;
	6525 : 1;
	6526 : 1;
	6527 : 1;
	6528 : 1;
	6529 : 1;
	6530 : 1;
	6531 : 1;
	6532 : 1;
	6533 : 1;
	6534 : 1;
	6535 : 1;
	6536 : 1;
	6537 : 1;
	6538 : 1;
	6539 : 1;
	6540 : 1;
	6541 : 1;
	6542 : 1;
	6543 : 1;
	6544 : 1;
	6545 : 1;
	6546 : 1;
	6547 : 1;
	6548 : 1;
	6549 : 1;
	6550 : 1;
	6551 : 1;
	6552 : 1;
	6553 : 1;
	6554 : 1;
	6555 : 1;
	6556 : 1;
	6557 : 1;
	6558 : 1;
	6559 : 1;
	6560 : 1;
	6561 : 1;
	6562 : 1;
	6563 : 1;
	6564 : 1;
	6565 : 1;
	6566 : 1;
	6567 : 1;
	6568 : 1;
	6569 : 1;
	6570 : 1;
	6571 : 1;
	6572 : 1;
	6573 : 1;
	6574 : 1;
	6575 : 1;
	6576 : 1;
	6577 : 1;
	6578 : 1;
	6579 : 1;
	6580 : 1;
	6581 : 1;
	6582 : 1;
	6583 : 1;
	6584 : 1;
	6585 : 1;
	6586 : 1;
	6587 : 1;
	6588 : 1;
	6589 : 1;
	6590 : 1;
	6591 : 1;
	6592 : 1;
	6593 : 1;
	6594 : 1;
	6595 : 1;
	6596 : 1;
	6597 : 1;
	6598 : 1;
	6599 : 1;
	6600 : 1;
	6601 : 1;
	6602 : 1;
	6603 : 1;
	6604 : 1;
	6605 : 1;
	6606 : 1;
	6607 : 1;
	6608 : 1;
	6609 : 1;
	6610 : 1;
	6611 : 1;
	6612 : 1;
	6613 : 1;
	6614 : 1;
	6615 : 1;
	6616 : 1;
	6617 : 1;
	6618 : 1;
	6619 : 1;
	6620 : 1;
	6621 : 1;
	6622 : 1;
	6623 : 1;
	6624 : 1;
	6625 : 1;
	6626 : 1;
	6627 : 1;
	6628 : 1;
	6629 : 1;
	6630 : 1;
	6631 : 1;
	6632 : 1;
	6633 : 1;
	6634 : 1;
	6635 : 1;
	6636 : 1;
	6637 : 1;
	6638 : 1;
	6639 : 1;
	6640 : 1;
	6641 : 1;
	6642 : 1;
	6643 : 1;
	6644 : 1;
	6645 : 1;
	6646 : 1;
	6647 : 1;
	6648 : 1;
	6649 : 1;
	6650 : 1;
	6651 : 1;
	6652 : 1;
	6653 : 1;
	6654 : 1;
	6655 : 1;
	6656 : 1;
	6657 : 1;
	6658 : 1;
	6659 : 1;
	6660 : 1;
	6661 : 1;
	6662 : 1;
	6663 : 1;
	6664 : 1;
	6665 : 1;
	6666 : 1;
	6667 : 1;
	6668 : 1;
	6669 : 1;
	6670 : 1;
	6671 : 1;
	6672 : 1;
	6673 : 1;
	6674 : 1;
	6675 : 1;
	6676 : 1;
	6677 : 1;
	6678 : 1;
	6679 : 1;
	6680 : 1;
	6681 : 1;
	6682 : 1;
	6683 : 1;
	6684 : 1;
	6685 : 1;
	6686 : 1;
	6687 : 1;
	6688 : 1;
	6689 : 1;
	6690 : 1;
	6691 : 1;
	6692 : 1;
	6693 : 1;
	6694 : 1;
	6695 : 1;
	6696 : 1;
	6697 : 1;
	6698 : 1;
	6699 : 1;
	6700 : 1;
	6701 : 1;
	6702 : 1;
	6703 : 1;
	6704 : 1;
	6705 : 1;
	6706 : 1;
	6707 : 1;
	6708 : 1;
	6709 : 1;
	6710 : 1;
	6711 : 1;
	6712 : 1;
	6713 : 1;
	6714 : 1;
	6715 : 1;
	6716 : 1;
	6717 : 1;
	6718 : 1;
	6719 : 1;
	6720 : 1;
	6721 : 1;
	6722 : 1;
	6723 : 1;
	6724 : 1;
	6725 : 1;
	6726 : 1;
	6727 : 1;
	6728 : 1;
	6729 : 1;
	6730 : 1;
	6731 : 1;
	6732 : 1;
	6733 : 1;
	6734 : 1;
	6735 : 1;
	6736 : 1;
	6737 : 1;
	6738 : 1;
	6739 : 1;
	6740 : 1;
	6741 : 1;
	6742 : 1;
	6743 : 1;
	6744 : 1;
	6745 : 1;
	6746 : 1;
	6747 : 1;
	6748 : 1;
	6749 : 1;
	6750 : 1;
	6751 : 1;
	6752 : 1;
	6753 : 1;
	6754 : 1;
	6755 : 1;
	6756 : 1;
	6757 : 1;
	6758 : 1;
	6759 : 1;
	6760 : 1;
	6761 : 1;
	6762 : 1;
	6763 : 1;
	6764 : 1;
	6765 : 1;
	6766 : 1;
	6767 : 1;
	6768 : 1;
	6769 : 1;
	6770 : 1;
	6771 : 1;
	6772 : 1;
	6773 : 1;
	6774 : 1;
	6775 : 1;
	6776 : 1;
	6777 : 1;
	6778 : 1;
	6779 : 1;
	6780 : 1;
	6781 : 1;
	6782 : 1;
	6783 : 1;
	6784 : 1;
	6785 : 1;
	6786 : 1;
	6787 : 1;
	6788 : 1;
	6789 : 1;
	6790 : 1;
	6791 : 1;
	6792 : 1;
	6793 : 1;
	6794 : 1;
	6795 : 1;
	6796 : 1;
	6797 : 1;
	6798 : 1;
	6799 : 1;
	6800 : 1;
	6801 : 1;
	6802 : 1;
	6803 : 1;
	6804 : 1;
	6805 : 1;
	6806 : 1;
	6807 : 1;
	6808 : 1;
	6809 : 1;
	6810 : 1;
	6811 : 1;
	6812 : 1;
	6813 : 1;
	6814 : 1;
	6815 : 1;
	6816 : 1;
	6817 : 1;
	6818 : 1;
	6819 : 1;
	6820 : 1;
	6821 : 1;
	6822 : 1;
	6823 : 1;
	6824 : 1;
	6825 : 1;
	6826 : 1;
	6827 : 1;
	6828 : 1;
	6829 : 1;
	6830 : 1;
	6831 : 1;
	6832 : 1;
	6833 : 1;
	6834 : 1;
	6835 : 1;
	6836 : 1;
	6837 : 1;
	6838 : 1;
	6839 : 1;
	6840 : 1;
	6841 : 1;
	6842 : 1;
	6843 : 1;
	6844 : 1;
	6845 : 1;
	6846 : 1;
	6847 : 1;
	6848 : 1;
	6849 : 1;
	6850 : 1;
	6851 : 1;
	6852 : 1;
	6853 : 1;
	6854 : 1;
	6855 : 1;
	6856 : 1;
	6857 : 1;
	6858 : 1;
	6859 : 1;
	6860 : 1;
	6861 : 1;
	6862 : 1;
	6863 : 1;
	6864 : 1;
	6865 : 1;
	6866 : 1;
	6867 : 1;
	6868 : 1;
	6869 : 1;
	6870 : 1;
	6871 : 1;
	6872 : 1;
	6873 : 1;
	6874 : 1;
	6875 : 1;
	6876 : 1;
	6877 : 1;
	6878 : 1;
	6879 : 1;
	6880 : 1;
	6881 : 1;
	6882 : 1;
	6883 : 1;
	6884 : 1;
	6885 : 1;
	6886 : 1;
	6887 : 1;
	6888 : 1;
	6889 : 1;
	6890 : 0;
	6891 : 1;
	6892 : 1;
	6893 : 0;
	6894 : 1;
	6895 : 1;
	6896 : 1;
	6897 : 1;
	6898 : 1;
	6899 : 1;
	6900 : 1;
	6901 : 0;
	6902 : 1;
	6903 : 1;
	6904 : 1;
	6905 : 1;
	6906 : 1;
	6907 : 1;
	6908 : 1;
	6909 : 1;
	6910 : 1;
	6911 : 1;
	6912 : 1;
	6913 : 1;
	6914 : 1;
	6915 : 1;
	6916 : 1;
	6917 : 1;
	6918 : 1;
	6919 : 1;
	6920 : 1;
	6921 : 1;
	6922 : 1;
	6923 : 1;
	6924 : 1;
	6925 : 1;
	6926 : 1;
	6927 : 1;
	6928 : 1;
	6929 : 1;
	6930 : 1;
	6931 : 1;
	6932 : 1;
	6933 : 1;
	6934 : 1;
	6935 : 1;
	6936 : 1;
	6937 : 1;
	6938 : 1;
	6939 : 1;
	6940 : 1;
	6941 : 1;
	6942 : 1;
	6943 : 1;
	6944 : 1;
	6945 : 1;
	6946 : 1;
	6947 : 1;
	6948 : 1;
	6949 : 1;
	6950 : 1;
	6951 : 1;
	6952 : 1;
	6953 : 1;
	6954 : 1;
	6955 : 1;
	6956 : 1;
	6957 : 1;
	6958 : 1;
	6959 : 1;
	6960 : 1;
	6961 : 1;
	6962 : 1;
	6963 : 1;
	6964 : 1;
	6965 : 1;
	6966 : 1;
	6967 : 1;
	6968 : 1;
	6969 : 1;
	6970 : 1;
	6971 : 1;
	6972 : 1;
	6973 : 1;
	6974 : 1;
	6975 : 1;
	6976 : 1;
	6977 : 1;
	6978 : 1;
	6979 : 1;
	6980 : 1;
	6981 : 1;
	6982 : 1;
	6983 : 1;
	6984 : 1;
	6985 : 1;
	6986 : 1;
	6987 : 1;
	6988 : 1;
	6989 : 1;
	6990 : 1;
	6991 : 1;
	6992 : 1;
	6993 : 1;
	6994 : 1;
	6995 : 1;
	6996 : 1;
	6997 : 1;
	6998 : 1;
	6999 : 1;
	7000 : 1;
	7001 : 1;
	7002 : 1;
	7003 : 1;
	7004 : 1;
	7005 : 1;
	7006 : 1;
	7007 : 1;
	7008 : 1;
	7009 : 1;
	7010 : 1;
	7011 : 1;
	7012 : 1;
	7013 : 1;
	7014 : 1;
	7015 : 1;
	7016 : 1;
	7017 : 1;
	7018 : 1;
	7019 : 1;
	7020 : 1;
	7021 : 1;
	7022 : 1;
	7023 : 1;
	7024 : 1;
	7025 : 1;
	7026 : 1;
	7027 : 1;
	7028 : 1;
	7029 : 1;
	7030 : 1;
	7031 : 1;
	7032 : 1;
	7033 : 1;
	7034 : 1;
	7035 : 1;
	7036 : 1;
	7037 : 1;
	7038 : 1;
	7039 : 1;
	7040 : 1;
	7041 : 1;
	7042 : 1;
	7043 : 1;
	7044 : 1;
	7045 : 1;
	7046 : 1;
	7047 : 1;
	7048 : 1;
	7049 : 1;
	7050 : 1;
	7051 : 1;
	7052 : 1;
	7053 : 1;
	7054 : 1;
	7055 : 1;
	7056 : 1;
	7057 : 1;
	7058 : 1;
	7059 : 1;
	7060 : 1;
	7061 : 1;
	7062 : 1;
	7063 : 1;
	7064 : 1;
	7065 : 1;
	7066 : 1;
	7067 : 1;
	7068 : 1;
	7069 : 1;
	7070 : 1;
	7071 : 1;
	7072 : 1;
	7073 : 1;
	7074 : 1;
	7075 : 1;
	7076 : 1;
	7077 : 1;
	7078 : 1;
	7079 : 1;
	7080 : 1;
	7081 : 1;
	7082 : 1;
	7083 : 1;
	7084 : 1;
	7085 : 1;
	7086 : 1;
	7087 : 1;
	7088 : 1;
	7089 : 1;
	7090 : 1;
	7091 : 1;
	7092 : 1;
	7093 : 1;
	7094 : 1;
	7095 : 1;
	7096 : 1;
	7097 : 1;
	7098 : 1;
	7099 : 1;
	7100 : 1;
	7101 : 1;
	7102 : 1;
	7103 : 1;
	7104 : 1;
	7105 : 1;
	7106 : 1;
	7107 : 1;
	7108 : 1;
	7109 : 1;
	7110 : 1;
	7111 : 1;
	7112 : 1;
	7113 : 1;
	7114 : 1;
	7115 : 1;
	7116 : 1;
	7117 : 1;
	7118 : 1;
	7119 : 1;
	7120 : 1;
	7121 : 1;
	7122 : 1;
	7123 : 1;
	7124 : 1;
	7125 : 1;
	7126 : 1;
	7127 : 1;
	7128 : 1;
	7129 : 0;
	7130 : 0;
	7131 : 0;
	7132 : 0;
	7133 : 0;
	7134 : 0;
	7135 : 1;
	7136 : 1;
	7137 : 1;
	7138 : 1;
	7139 : 1;
	7140 : 1;
	7141 : 0;
	7142 : 0;
	7143 : 1;
	7144 : 1;
	7145 : 1;
	7146 : 1;
	7147 : 1;
	7148 : 1;
	7149 : 1;
	7150 : 1;
	7151 : 1;
	7152 : 1;
	7153 : 1;
	7154 : 1;
	7155 : 1;
	7156 : 1;
	7157 : 1;
	7158 : 1;
	7159 : 1;
	7160 : 1;
	7161 : 1;
	7162 : 1;
	7163 : 1;
	7164 : 1;
	7165 : 1;
	7166 : 1;
	7167 : 1;
	7168 : 1;
	7169 : 1;
	7170 : 1;
	7171 : 1;
	7172 : 1;
	7173 : 1;
	7174 : 1;
	7175 : 1;
	7176 : 1;
	7177 : 1;
	7178 : 1;
	7179 : 1;
	7180 : 1;
	7181 : 1;
	7182 : 1;
	7183 : 1;
	7184 : 1;
	7185 : 1;
	7186 : 1;
	7187 : 1;
	7188 : 1;
	7189 : 1;
	7190 : 1;
	7191 : 1;
	7192 : 1;
	7193 : 1;
	7194 : 1;
	7195 : 1;
	7196 : 1;
	7197 : 1;
	7198 : 1;
	7199 : 1;
	7200 : 1;
	7201 : 1;
	7202 : 1;
	7203 : 1;
	7204 : 1;
	7205 : 1;
	7206 : 1;
	7207 : 1;
	7208 : 1;
	7209 : 1;
	7210 : 1;
	7211 : 1;
	7212 : 1;
	7213 : 1;
	7214 : 1;
	7215 : 1;
	7216 : 1;
	7217 : 1;
	7218 : 1;
	7219 : 1;
	7220 : 1;
	7221 : 1;
	7222 : 1;
	7223 : 1;
	7224 : 1;
	7225 : 1;
	7226 : 1;
	7227 : 1;
	7228 : 1;
	7229 : 1;
	7230 : 1;
	7231 : 1;
	7232 : 1;
	7233 : 1;
	7234 : 1;
	7235 : 1;
	7236 : 1;
	7237 : 1;
	7238 : 1;
	7239 : 1;
	7240 : 1;
	7241 : 1;
	7242 : 1;
	7243 : 1;
	7244 : 1;
	7245 : 1;
	7246 : 1;
	7247 : 1;
	7248 : 1;
	7249 : 1;
	7250 : 1;
	7251 : 1;
	7252 : 1;
	7253 : 1;
	7254 : 1;
	7255 : 1;
	7256 : 1;
	7257 : 1;
	7258 : 1;
	7259 : 1;
	7260 : 1;
	7261 : 1;
	7262 : 1;
	7263 : 1;
	7264 : 1;
	7265 : 1;
	7266 : 1;
	7267 : 1;
	7268 : 1;
	7269 : 1;
	7270 : 1;
	7271 : 1;
	7272 : 1;
	7273 : 1;
	7274 : 1;
	7275 : 1;
	7276 : 1;
	7277 : 1;
	7278 : 1;
	7279 : 1;
	7280 : 1;
	7281 : 1;
	7282 : 1;
	7283 : 1;
	7284 : 1;
	7285 : 1;
	7286 : 1;
	7287 : 1;
	7288 : 1;
	7289 : 1;
	7290 : 1;
	7291 : 1;
	7292 : 1;
	7293 : 1;
	7294 : 1;
	7295 : 1;
	7296 : 1;
	7297 : 1;
	7298 : 1;
	7299 : 1;
	7300 : 1;
	7301 : 1;
	7302 : 1;
	7303 : 1;
	7304 : 1;
	7305 : 1;
	7306 : 1;
	7307 : 1;
	7308 : 1;
	7309 : 1;
	7310 : 1;
	7311 : 1;
	7312 : 1;
	7313 : 1;
	7314 : 1;
	7315 : 1;
	7316 : 1;
	7317 : 1;
	7318 : 1;
	7319 : 1;
	7320 : 1;
	7321 : 1;
	7322 : 1;
	7323 : 1;
	7324 : 1;
	7325 : 1;
	7326 : 1;
	7327 : 1;
	7328 : 1;
	7329 : 1;
	7330 : 1;
	7331 : 1;
	7332 : 1;
	7333 : 1;
	7334 : 1;
	7335 : 1;
	7336 : 1;
	7337 : 1;
	7338 : 1;
	7339 : 1;
	7340 : 1;
	7341 : 1;
	7342 : 1;
	7343 : 1;
	7344 : 1;
	7345 : 1;
	7346 : 1;
	7347 : 1;
	7348 : 1;
	7349 : 1;
	7350 : 1;
	7351 : 1;
	7352 : 1;
	7353 : 1;
	7354 : 1;
	7355 : 1;
	7356 : 1;
	7357 : 1;
	7358 : 1;
	7359 : 1;
	7360 : 1;
	7361 : 1;
	7362 : 1;
	7363 : 1;
	7364 : 1;
	7365 : 1;
	7366 : 1;
	7367 : 1;
	7368 : 1;
	7369 : 1;
	7370 : 0;
	7371 : 0;
	7372 : 1;
	7373 : 0;
	7374 : 0;
	7375 : 1;
	7376 : 1;
	7377 : 1;
	7378 : 1;
	7379 : 1;
	7380 : 1;
	7381 : 1;
	7382 : 0;
	7383 : 1;
	7384 : 1;
	7385 : 1;
	7386 : 1;
	7387 : 1;
	7388 : 1;
	7389 : 1;
	7390 : 1;
	7391 : 1;
	7392 : 1;
	7393 : 1;
	7394 : 1;
	7395 : 1;
	7396 : 1;
	7397 : 1;
	7398 : 1;
	7399 : 1;
	7400 : 1;
	7401 : 1;
	7402 : 1;
	7403 : 1;
	7404 : 1;
	7405 : 1;
	7406 : 1;
	7407 : 1;
	7408 : 1;
	7409 : 1;
	7410 : 1;
	7411 : 1;
	7412 : 1;
	7413 : 1;
	7414 : 1;
	7415 : 1;
	7416 : 1;
	7417 : 1;
	7418 : 1;
	7419 : 1;
	7420 : 1;
	7421 : 1;
	7422 : 1;
	7423 : 1;
	7424 : 1;
	7425 : 1;
	7426 : 1;
	7427 : 1;
	7428 : 1;
	7429 : 1;
	7430 : 1;
	7431 : 1;
	7432 : 1;
	7433 : 1;
	7434 : 1;
	7435 : 1;
	7436 : 1;
	7437 : 1;
	7438 : 1;
	7439 : 1;
	7440 : 1;
	7441 : 1;
	7442 : 1;
	7443 : 1;
	7444 : 1;
	7445 : 1;
	7446 : 1;
	7447 : 1;
	7448 : 1;
	7449 : 1;
	7450 : 1;
	7451 : 1;
	7452 : 1;
	7453 : 1;
	7454 : 1;
	7455 : 1;
	7456 : 1;
	7457 : 1;
	7458 : 1;
	7459 : 1;
	7460 : 1;
	7461 : 1;
	7462 : 1;
	7463 : 1;
	7464 : 1;
	7465 : 1;
	7466 : 1;
	7467 : 1;
	7468 : 1;
	7469 : 1;
	7470 : 1;
	7471 : 1;
	7472 : 1;
	7473 : 1;
	7474 : 1;
	7475 : 1;
	7476 : 1;
	7477 : 1;
	7478 : 1;
	7479 : 1;
	7480 : 1;
	7481 : 1;
	7482 : 1;
	7483 : 1;
	7484 : 1;
	7485 : 1;
	7486 : 1;
	7487 : 1;
	7488 : 1;
	7489 : 1;
	7490 : 1;
	7491 : 1;
	7492 : 1;
	7493 : 1;
	7494 : 1;
	7495 : 1;
	7496 : 1;
	7497 : 1;
	7498 : 1;
	7499 : 1;
	7500 : 1;
	7501 : 1;
	7502 : 1;
	7503 : 1;
	7504 : 1;
	7505 : 1;
	7506 : 1;
	7507 : 1;
	7508 : 1;
	7509 : 1;
	7510 : 1;
	7511 : 1;
	7512 : 1;
	7513 : 1;
	7514 : 1;
	7515 : 1;
	7516 : 1;
	7517 : 1;
	7518 : 1;
	7519 : 1;
	7520 : 1;
	7521 : 1;
	7522 : 1;
	7523 : 1;
	7524 : 1;
	7525 : 1;
	7526 : 1;
	7527 : 1;
	7528 : 1;
	7529 : 1;
	7530 : 1;
	7531 : 1;
	7532 : 1;
	7533 : 1;
	7534 : 1;
	7535 : 1;
	7536 : 1;
	7537 : 1;
	7538 : 1;
	7539 : 1;
	7540 : 1;
	7541 : 1;
	7542 : 1;
	7543 : 1;
	7544 : 1;
	7545 : 1;
	7546 : 1;
	7547 : 1;
	7548 : 1;
	7549 : 1;
	7550 : 1;
	7551 : 1;
	7552 : 1;
	7553 : 1;
	7554 : 1;
	7555 : 1;
	7556 : 1;
	7557 : 1;
	7558 : 1;
	7559 : 1;
	7560 : 1;
	7561 : 1;
	7562 : 1;
	7563 : 1;
	7564 : 1;
	7565 : 1;
	7566 : 1;
	7567 : 1;
	7568 : 1;
	7569 : 1;
	7570 : 1;
	7571 : 1;
	7572 : 1;
	7573 : 1;
	7574 : 1;
	7575 : 1;
	7576 : 1;
	7577 : 1;
	7578 : 1;
	7579 : 1;
	7580 : 1;
	7581 : 1;
	7582 : 1;
	7583 : 1;
	7584 : 1;
	7585 : 1;
	7586 : 1;
	7587 : 1;
	7588 : 1;
	7589 : 1;
	7590 : 1;
	7591 : 1;
	7592 : 1;
	7593 : 1;
	7594 : 1;
	7595 : 1;
	7596 : 1;
	7597 : 1;
	7598 : 1;
	7599 : 1;
	7600 : 1;
	7601 : 1;
	7602 : 1;
	7603 : 1;
	7604 : 1;
	7605 : 1;
	7606 : 1;
	7607 : 0;
	7608 : 0;
	7609 : 1;
	7610 : 0;
	7611 : 1;
	7612 : 1;
	7613 : 0;
	7614 : 0;
	7615 : 1;
	7616 : 1;
	7617 : 1;
	7618 : 1;
	7619 : 1;
	7620 : 1;
	7621 : 1;
	7622 : 0;
	7623 : 1;
	7624 : 1;
	7625 : 1;
	7626 : 1;
	7627 : 1;
	7628 : 1;
	7629 : 1;
	7630 : 1;
	7631 : 1;
	7632 : 1;
	7633 : 1;
	7634 : 1;
	7635 : 1;
	7636 : 1;
	7637 : 1;
	7638 : 1;
	7639 : 1;
	7640 : 1;
	7641 : 1;
	7642 : 1;
	7643 : 1;
	7644 : 1;
	7645 : 1;
	7646 : 1;
	7647 : 1;
	7648 : 1;
	7649 : 1;
	7650 : 1;
	7651 : 1;
	7652 : 1;
	7653 : 1;
	7654 : 1;
	7655 : 1;
	7656 : 1;
	7657 : 1;
	7658 : 1;
	7659 : 1;
	7660 : 1;
	7661 : 1;
	7662 : 1;
	7663 : 1;
	7664 : 1;
	7665 : 1;
	7666 : 1;
	7667 : 1;
	7668 : 1;
	7669 : 1;
	7670 : 1;
	7671 : 1;
	7672 : 1;
	7673 : 1;
	7674 : 1;
	7675 : 1;
	7676 : 1;
	7677 : 1;
	7678 : 1;
	7679 : 1;
	7680 : 1;
	7681 : 1;
	7682 : 1;
	7683 : 1;
	7684 : 1;
	7685 : 1;
	7686 : 1;
	7687 : 1;
	7688 : 1;
	7689 : 1;
	7690 : 1;
	7691 : 1;
	7692 : 1;
	7693 : 1;
	7694 : 1;
	7695 : 1;
	7696 : 1;
	7697 : 1;
	7698 : 1;
	7699 : 1;
	7700 : 1;
	7701 : 1;
	7702 : 1;
	7703 : 1;
	7704 : 1;
	7705 : 1;
	7706 : 1;
	7707 : 1;
	7708 : 1;
	7709 : 1;
	7710 : 1;
	7711 : 1;
	7712 : 1;
	7713 : 1;
	7714 : 1;
	7715 : 1;
	7716 : 1;
	7717 : 1;
	7718 : 1;
	7719 : 1;
	7720 : 1;
	7721 : 1;
	7722 : 1;
	7723 : 1;
	7724 : 1;
	7725 : 1;
	7726 : 1;
	7727 : 1;
	7728 : 1;
	7729 : 1;
	7730 : 1;
	7731 : 1;
	7732 : 1;
	7733 : 1;
	7734 : 1;
	7735 : 1;
	7736 : 1;
	7737 : 1;
	7738 : 1;
	7739 : 1;
	7740 : 1;
	7741 : 1;
	7742 : 1;
	7743 : 1;
	7744 : 1;
	7745 : 1;
	7746 : 1;
	7747 : 1;
	7748 : 1;
	7749 : 1;
	7750 : 1;
	7751 : 1;
	7752 : 1;
	7753 : 1;
	7754 : 1;
	7755 : 1;
	7756 : 1;
	7757 : 1;
	7758 : 1;
	7759 : 1;
	7760 : 1;
	7761 : 1;
	7762 : 1;
	7763 : 1;
	7764 : 1;
	7765 : 1;
	7766 : 1;
	7767 : 1;
	7768 : 1;
	7769 : 1;
	7770 : 1;
	7771 : 1;
	7772 : 1;
	7773 : 1;
	7774 : 1;
	7775 : 1;
	7776 : 1;
	7777 : 1;
	7778 : 1;
	7779 : 1;
	7780 : 1;
	7781 : 1;
	7782 : 1;
	7783 : 1;
	7784 : 1;
	7785 : 1;
	7786 : 1;
	7787 : 1;
	7788 : 1;
	7789 : 1;
	7790 : 1;
	7791 : 1;
	7792 : 1;
	7793 : 1;
	7794 : 1;
	7795 : 1;
	7796 : 1;
	7797 : 1;
	7798 : 1;
	7799 : 1;
	7800 : 1;
	7801 : 1;
	7802 : 1;
	7803 : 1;
	7804 : 1;
	7805 : 1;
	7806 : 1;
	7807 : 1;
	7808 : 1;
	7809 : 1;
	7810 : 1;
	7811 : 1;
	7812 : 1;
	7813 : 1;
	7814 : 1;
	7815 : 1;
	7816 : 1;
	7817 : 1;
	7818 : 1;
	7819 : 1;
	7820 : 1;
	7821 : 1;
	7822 : 1;
	7823 : 1;
	7824 : 1;
	7825 : 1;
	7826 : 1;
	7827 : 1;
	7828 : 1;
	7829 : 1;
	7830 : 1;
	7831 : 1;
	7832 : 1;
	7833 : 1;
	7834 : 1;
	7835 : 1;
	7836 : 1;
	7837 : 1;
	7838 : 1;
	7839 : 1;
	7840 : 1;
	7841 : 1;
	7842 : 1;
	7843 : 1;
	7844 : 1;
	7845 : 1;
	7846 : 1;
	7847 : 0;
	7848 : 0;
	7849 : 1;
	7850 : 1;
	7851 : 1;
	7852 : 1;
	7853 : 0;
	7854 : 1;
	7855 : 1;
	7856 : 1;
	7857 : 1;
	7858 : 1;
	7859 : 1;
	7860 : 1;
	7861 : 1;
	7862 : 0;
	7863 : 1;
	7864 : 1;
	7865 : 1;
	7866 : 1;
	7867 : 1;
	7868 : 1;
	7869 : 1;
	7870 : 1;
	7871 : 1;
	7872 : 1;
	7873 : 1;
	7874 : 1;
	7875 : 1;
	7876 : 1;
	7877 : 1;
	7878 : 1;
	7879 : 1;
	7880 : 1;
	7881 : 1;
	7882 : 1;
	7883 : 1;
	7884 : 1;
	7885 : 1;
	7886 : 1;
	7887 : 1;
	7888 : 1;
	7889 : 1;
	7890 : 1;
	7891 : 1;
	7892 : 1;
	7893 : 1;
	7894 : 1;
	7895 : 1;
	7896 : 1;
	7897 : 1;
	7898 : 1;
	7899 : 1;
	7900 : 1;
	7901 : 1;
	7902 : 1;
	7903 : 1;
	7904 : 1;
	7905 : 1;
	7906 : 1;
	7907 : 1;
	7908 : 1;
	7909 : 1;
	7910 : 1;
	7911 : 1;
	7912 : 1;
	7913 : 1;
	7914 : 1;
	7915 : 1;
	7916 : 1;
	7917 : 1;
	7918 : 1;
	7919 : 1;
	7920 : 1;
	7921 : 1;
	7922 : 1;
	7923 : 1;
	7924 : 1;
	7925 : 1;
	7926 : 1;
	7927 : 1;
	7928 : 1;
	7929 : 1;
	7930 : 1;
	7931 : 1;
	7932 : 1;
	7933 : 1;
	7934 : 1;
	7935 : 1;
	7936 : 1;
	7937 : 1;
	7938 : 1;
	7939 : 1;
	7940 : 1;
	7941 : 1;
	7942 : 1;
	7943 : 1;
	7944 : 1;
	7945 : 1;
	7946 : 1;
	7947 : 1;
	7948 : 1;
	7949 : 1;
	7950 : 1;
	7951 : 1;
	7952 : 1;
	7953 : 1;
	7954 : 1;
	7955 : 1;
	7956 : 1;
	7957 : 1;
	7958 : 1;
	7959 : 1;
	7960 : 1;
	7961 : 1;
	7962 : 1;
	7963 : 1;
	7964 : 1;
	7965 : 1;
	7966 : 1;
	7967 : 1;
	7968 : 1;
	7969 : 1;
	7970 : 1;
	7971 : 1;
	7972 : 1;
	7973 : 1;
	7974 : 1;
	7975 : 1;
	7976 : 1;
	7977 : 1;
	7978 : 1;
	7979 : 1;
	7980 : 1;
	7981 : 1;
	7982 : 1;
	7983 : 1;
	7984 : 1;
	7985 : 1;
	7986 : 1;
	7987 : 1;
	7988 : 1;
	7989 : 1;
	7990 : 1;
	7991 : 1;
	7992 : 0;
	7993 : 1;
	7994 : 1;
	7995 : 1;
	7996 : 1;
	7997 : 1;
	7998 : 1;
	7999 : 1;
	8000 : 1;
	8001 : 1;
	8002 : 1;
	8003 : 1;
	8004 : 1;
	8005 : 1;
	8006 : 1;
	8007 : 1;
	8008 : 1;
	8009 : 1;
	8010 : 1;
	8011 : 1;
	8012 : 1;
	8013 : 1;
	8014 : 1;
	8015 : 1;
	8016 : 1;
	8017 : 1;
	8018 : 1;
	8019 : 1;
	8020 : 1;
	8021 : 1;
	8022 : 0;
	8023 : 0;
	8024 : 0;
	8025 : 0;
	8026 : 0;
	8027 : 1;
	8028 : 0;
	8029 : 1;
	8030 : 1;
	8031 : 1;
	8032 : 1;
	8033 : 1;
	8034 : 1;
	8035 : 1;
	8036 : 1;
	8037 : 1;
	8038 : 1;
	8039 : 1;
	8040 : 1;
	8041 : 1;
	8042 : 0;
	8043 : 0;
	8044 : 1;
	8045 : 1;
	8046 : 1;
	8047 : 0;
	8048 : 0;
	8049 : 0;
	8050 : 0;
	8051 : 1;
	8052 : 1;
	8053 : 1;
	8054 : 1;
	8055 : 1;
	8056 : 1;
	8057 : 1;
	8058 : 1;
	8059 : 1;
	8060 : 1;
	8061 : 1;
	8062 : 1;
	8063 : 1;
	8064 : 1;
	8065 : 1;
	8066 : 1;
	8067 : 1;
	8068 : 0;
	8069 : 1;
	8070 : 1;
	8071 : 1;
	8072 : 1;
	8073 : 1;
	8074 : 1;
	8075 : 1;
	8076 : 1;
	8077 : 1;
	8078 : 1;
	8079 : 1;
	8080 : 1;
	8081 : 1;
	8082 : 1;
	8083 : 1;
	8084 : 1;
	8085 : 1;
	8086 : 1;
	8087 : 0;
	8088 : 0;
	8089 : 1;
	8090 : 1;
	8091 : 1;
	8092 : 1;
	8093 : 1;
	8094 : 1;
	8095 : 1;
	8096 : 1;
	8097 : 1;
	8098 : 1;
	8099 : 1;
	8100 : 1;
	8101 : 1;
	8102 : 0;
	8103 : 1;
	8104 : 1;
	8105 : 1;
	8106 : 1;
	8107 : 1;
	8108 : 1;
	8109 : 1;
	8110 : 1;
	8111 : 1;
	8112 : 1;
	8113 : 1;
	8114 : 1;
	8115 : 1;
	8116 : 1;
	8117 : 1;
	8118 : 1;
	8119 : 1;
	8120 : 1;
	8121 : 1;
	8122 : 1;
	8123 : 1;
	8124 : 1;
	8125 : 1;
	8126 : 1;
	8127 : 1;
	8128 : 1;
	8129 : 1;
	8130 : 1;
	8131 : 1;
	8132 : 1;
	8133 : 1;
	8134 : 1;
	8135 : 1;
	8136 : 1;
	8137 : 1;
	8138 : 1;
	8139 : 1;
	8140 : 1;
	8141 : 1;
	8142 : 1;
	8143 : 1;
	8144 : 1;
	8145 : 1;
	8146 : 1;
	8147 : 1;
	8148 : 1;
	8149 : 1;
	8150 : 1;
	8151 : 1;
	8152 : 1;
	8153 : 1;
	8154 : 1;
	8155 : 1;
	8156 : 1;
	8157 : 1;
	8158 : 1;
	8159 : 1;
	8160 : 1;
	8161 : 1;
	8162 : 1;
	8163 : 1;
	8164 : 1;
	8165 : 1;
	8166 : 1;
	8167 : 1;
	8168 : 1;
	8169 : 1;
	8170 : 1;
	8171 : 1;
	8172 : 1;
	8173 : 1;
	8174 : 1;
	8175 : 1;
	8176 : 1;
	8177 : 1;
	8178 : 1;
	8179 : 1;
	8180 : 1;
	8181 : 1;
	8182 : 1;
	8183 : 1;
	8184 : 1;
	8185 : 1;
	8186 : 1;
	8187 : 1;
	8188 : 1;
	8189 : 1;
	8190 : 1;
	8191 : 1;
	8192 : 1;
	8193 : 1;
	8194 : 1;
	8195 : 1;
	8196 : 1;
	8197 : 1;
	8198 : 1;
	8199 : 1;
	8200 : 1;
	8201 : 1;
	8202 : 1;
	8203 : 1;
	8204 : 1;
	8205 : 1;
	8206 : 1;
	8207 : 1;
	8208 : 1;
	8209 : 1;
	8210 : 1;
	8211 : 1;
	8212 : 1;
	8213 : 1;
	8214 : 1;
	8215 : 1;
	8216 : 1;
	8217 : 1;
	8218 : 1;
	8219 : 1;
	8220 : 1;
	8221 : 1;
	8222 : 1;
	8223 : 1;
	8224 : 1;
	8225 : 1;
	8226 : 1;
	8227 : 1;
	8228 : 1;
	8229 : 1;
	8230 : 1;
	8231 : 1;
	8232 : 0;
	8233 : 1;
	8234 : 1;
	8235 : 1;
	8236 : 1;
	8237 : 1;
	8238 : 1;
	8239 : 1;
	8240 : 1;
	8241 : 1;
	8242 : 1;
	8243 : 1;
	8244 : 1;
	8245 : 1;
	8246 : 1;
	8247 : 1;
	8248 : 1;
	8249 : 1;
	8250 : 1;
	8251 : 1;
	8252 : 1;
	8253 : 1;
	8254 : 1;
	8255 : 1;
	8256 : 1;
	8257 : 1;
	8258 : 1;
	8259 : 1;
	8260 : 1;
	8261 : 1;
	8262 : 0;
	8263 : 1;
	8264 : 1;
	8265 : 1;
	8266 : 1;
	8267 : 1;
	8268 : 1;
	8269 : 1;
	8270 : 1;
	8271 : 1;
	8272 : 1;
	8273 : 1;
	8274 : 1;
	8275 : 1;
	8276 : 1;
	8277 : 1;
	8278 : 1;
	8279 : 1;
	8280 : 1;
	8281 : 1;
	8282 : 0;
	8283 : 0;
	8284 : 1;
	8285 : 1;
	8286 : 1;
	8287 : 0;
	8288 : 1;
	8289 : 1;
	8290 : 1;
	8291 : 0;
	8292 : 1;
	8293 : 1;
	8294 : 1;
	8295 : 1;
	8296 : 1;
	8297 : 1;
	8298 : 1;
	8299 : 1;
	8300 : 1;
	8301 : 1;
	8302 : 1;
	8303 : 1;
	8304 : 1;
	8305 : 1;
	8306 : 1;
	8307 : 1;
	8308 : 1;
	8309 : 1;
	8310 : 1;
	8311 : 1;
	8312 : 1;
	8313 : 1;
	8314 : 1;
	8315 : 1;
	8316 : 1;
	8317 : 1;
	8318 : 1;
	8319 : 1;
	8320 : 1;
	8321 : 1;
	8322 : 1;
	8323 : 0;
	8324 : 1;
	8325 : 1;
	8326 : 1;
	8327 : 0;
	8328 : 0;
	8329 : 1;
	8330 : 1;
	8331 : 1;
	8332 : 1;
	8333 : 1;
	8334 : 1;
	8335 : 1;
	8336 : 1;
	8337 : 1;
	8338 : 0;
	8339 : 0;
	8340 : 1;
	8341 : 1;
	8342 : 0;
	8343 : 1;
	8344 : 1;
	8345 : 1;
	8346 : 1;
	8347 : 1;
	8348 : 1;
	8349 : 1;
	8350 : 1;
	8351 : 1;
	8352 : 1;
	8353 : 1;
	8354 : 1;
	8355 : 1;
	8356 : 1;
	8357 : 1;
	8358 : 1;
	8359 : 1;
	8360 : 1;
	8361 : 1;
	8362 : 1;
	8363 : 1;
	8364 : 1;
	8365 : 1;
	8366 : 1;
	8367 : 1;
	8368 : 1;
	8369 : 1;
	8370 : 1;
	8371 : 1;
	8372 : 1;
	8373 : 1;
	8374 : 1;
	8375 : 1;
	8376 : 1;
	8377 : 1;
	8378 : 1;
	8379 : 1;
	8380 : 1;
	8381 : 1;
	8382 : 1;
	8383 : 1;
	8384 : 1;
	8385 : 1;
	8386 : 1;
	8387 : 1;
	8388 : 1;
	8389 : 1;
	8390 : 1;
	8391 : 1;
	8392 : 1;
	8393 : 1;
	8394 : 1;
	8395 : 1;
	8396 : 1;
	8397 : 1;
	8398 : 1;
	8399 : 1;
	8400 : 1;
	8401 : 1;
	8402 : 1;
	8403 : 1;
	8404 : 1;
	8405 : 1;
	8406 : 1;
	8407 : 1;
	8408 : 1;
	8409 : 1;
	8410 : 1;
	8411 : 1;
	8412 : 1;
	8413 : 1;
	8414 : 1;
	8415 : 1;
	8416 : 1;
	8417 : 1;
	8418 : 1;
	8419 : 1;
	8420 : 1;
	8421 : 1;
	8422 : 1;
	8423 : 1;
	8424 : 1;
	8425 : 1;
	8426 : 1;
	8427 : 1;
	8428 : 1;
	8429 : 1;
	8430 : 1;
	8431 : 1;
	8432 : 1;
	8433 : 1;
	8434 : 1;
	8435 : 1;
	8436 : 1;
	8437 : 1;
	8438 : 1;
	8439 : 1;
	8440 : 1;
	8441 : 1;
	8442 : 1;
	8443 : 1;
	8444 : 1;
	8445 : 1;
	8446 : 1;
	8447 : 1;
	8448 : 1;
	8449 : 1;
	8450 : 1;
	8451 : 1;
	8452 : 1;
	8453 : 1;
	8454 : 1;
	8455 : 1;
	8456 : 1;
	8457 : 1;
	8458 : 1;
	8459 : 1;
	8460 : 1;
	8461 : 1;
	8462 : 1;
	8463 : 1;
	8464 : 1;
	8465 : 1;
	8466 : 1;
	8467 : 1;
	8468 : 1;
	8469 : 1;
	8470 : 1;
	8471 : 0;
	8472 : 0;
	8473 : 1;
	8474 : 1;
	8475 : 1;
	8476 : 1;
	8477 : 1;
	8478 : 1;
	8479 : 1;
	8480 : 1;
	8481 : 1;
	8482 : 1;
	8483 : 1;
	8484 : 1;
	8485 : 1;
	8486 : 1;
	8487 : 1;
	8488 : 1;
	8489 : 1;
	8490 : 1;
	8491 : 1;
	8492 : 1;
	8493 : 1;
	8494 : 1;
	8495 : 1;
	8496 : 1;
	8497 : 1;
	8498 : 1;
	8499 : 1;
	8500 : 1;
	8501 : 1;
	8502 : 0;
	8503 : 1;
	8504 : 1;
	8505 : 1;
	8506 : 1;
	8507 : 1;
	8508 : 1;
	8509 : 1;
	8510 : 1;
	8511 : 1;
	8512 : 1;
	8513 : 1;
	8514 : 1;
	8515 : 1;
	8516 : 1;
	8517 : 1;
	8518 : 1;
	8519 : 1;
	8520 : 1;
	8521 : 1;
	8522 : 0;
	8523 : 0;
	8524 : 1;
	8525 : 1;
	8526 : 1;
	8527 : 0;
	8528 : 1;
	8529 : 1;
	8530 : 1;
	8531 : 0;
	8532 : 1;
	8533 : 1;
	8534 : 1;
	8535 : 1;
	8536 : 1;
	8537 : 1;
	8538 : 1;
	8539 : 1;
	8540 : 1;
	8541 : 1;
	8542 : 1;
	8543 : 1;
	8544 : 1;
	8545 : 1;
	8546 : 1;
	8547 : 1;
	8548 : 1;
	8549 : 1;
	8550 : 1;
	8551 : 1;
	8552 : 1;
	8553 : 1;
	8554 : 1;
	8555 : 1;
	8556 : 1;
	8557 : 1;
	8558 : 1;
	8559 : 1;
	8560 : 1;
	8561 : 1;
	8562 : 1;
	8563 : 0;
	8564 : 0;
	8565 : 1;
	8566 : 1;
	8567 : 0;
	8568 : 0;
	8569 : 1;
	8570 : 1;
	8571 : 1;
	8572 : 1;
	8573 : 1;
	8574 : 1;
	8575 : 1;
	8576 : 1;
	8577 : 1;
	8578 : 0;
	8579 : 0;
	8580 : 1;
	8581 : 1;
	8582 : 0;
	8583 : 1;
	8584 : 1;
	8585 : 1;
	8586 : 1;
	8587 : 1;
	8588 : 1;
	8589 : 1;
	8590 : 1;
	8591 : 1;
	8592 : 1;
	8593 : 1;
	8594 : 1;
	8595 : 1;
	8596 : 1;
	8597 : 1;
	8598 : 1;
	8599 : 1;
	8600 : 1;
	8601 : 1;
	8602 : 1;
	8603 : 1;
	8604 : 1;
	8605 : 1;
	8606 : 1;
	8607 : 1;
	8608 : 1;
	8609 : 1;
	8610 : 1;
	8611 : 1;
	8612 : 1;
	8613 : 1;
	8614 : 1;
	8615 : 1;
	8616 : 1;
	8617 : 1;
	8618 : 1;
	8619 : 1;
	8620 : 1;
	8621 : 1;
	8622 : 1;
	8623 : 1;
	8624 : 1;
	8625 : 1;
	8626 : 1;
	8627 : 1;
	8628 : 1;
	8629 : 1;
	8630 : 1;
	8631 : 1;
	8632 : 1;
	8633 : 1;
	8634 : 1;
	8635 : 1;
	8636 : 1;
	8637 : 1;
	8638 : 1;
	8639 : 1;
	8640 : 1;
	8641 : 1;
	8642 : 1;
	8643 : 1;
	8644 : 1;
	8645 : 1;
	8646 : 1;
	8647 : 1;
	8648 : 1;
	8649 : 1;
	8650 : 1;
	8651 : 1;
	8652 : 1;
	8653 : 1;
	8654 : 1;
	8655 : 1;
	8656 : 1;
	8657 : 1;
	8658 : 1;
	8659 : 1;
	8660 : 1;
	8661 : 1;
	8662 : 1;
	8663 : 1;
	8664 : 1;
	8665 : 1;
	8666 : 1;
	8667 : 1;
	8668 : 1;
	8669 : 1;
	8670 : 1;
	8671 : 1;
	8672 : 1;
	8673 : 1;
	8674 : 1;
	8675 : 1;
	8676 : 1;
	8677 : 1;
	8678 : 1;
	8679 : 1;
	8680 : 1;
	8681 : 1;
	8682 : 1;
	8683 : 1;
	8684 : 1;
	8685 : 1;
	8686 : 1;
	8687 : 1;
	8688 : 1;
	8689 : 1;
	8690 : 1;
	8691 : 1;
	8692 : 1;
	8693 : 1;
	8694 : 1;
	8695 : 1;
	8696 : 1;
	8697 : 0;
	8698 : 0;
	8699 : 0;
	8700 : 0;
	8701 : 1;
	8702 : 0;
	8703 : 0;
	8704 : 0;
	8705 : 0;
	8706 : 1;
	8707 : 1;
	8708 : 0;
	8709 : 0;
	8710 : 0;
	8711 : 0;
	8712 : 0;
	8713 : 1;
	8714 : 1;
	8715 : 1;
	8716 : 0;
	8717 : 1;
	8718 : 1;
	8719 : 1;
	8720 : 0;
	8721 : 1;
	8722 : 1;
	8723 : 0;
	8724 : 0;
	8725 : 0;
	8726 : 0;
	8727 : 1;
	8728 : 0;
	8729 : 1;
	8730 : 1;
	8731 : 0;
	8732 : 0;
	8733 : 1;
	8734 : 0;
	8735 : 0;
	8736 : 0;
	8737 : 0;
	8738 : 0;
	8739 : 1;
	8740 : 1;
	8741 : 1;
	8742 : 0;
	8743 : 0;
	8744 : 0;
	8745 : 0;
	8746 : 1;
	8747 : 1;
	8748 : 0;
	8749 : 1;
	8750 : 0;
	8751 : 0;
	8752 : 0;
	8753 : 0;
	8754 : 1;
	8755 : 1;
	8756 : 0;
	8757 : 0;
	8758 : 0;
	8759 : 0;
	8760 : 0;
	8761 : 1;
	8762 : 0;
	8763 : 0;
	8764 : 1;
	8765 : 1;
	8766 : 1;
	8767 : 0;
	8768 : 1;
	8769 : 1;
	8770 : 1;
	8771 : 0;
	8772 : 1;
	8773 : 0;
	8774 : 1;
	8775 : 0;
	8776 : 0;
	8777 : 1;
	8778 : 1;
	8779 : 0;
	8780 : 0;
	8781 : 0;
	8782 : 0;
	8783 : 1;
	8784 : 1;
	8785 : 1;
	8786 : 1;
	8787 : 0;
	8788 : 0;
	8789 : 1;
	8790 : 0;
	8791 : 0;
	8792 : 0;
	8793 : 0;
	8794 : 1;
	8795 : 1;
	8796 : 1;
	8797 : 0;
	8798 : 0;
	8799 : 0;
	8800 : 0;
	8801 : 1;
	8802 : 0;
	8803 : 0;
	8804 : 0;
	8805 : 0;
	8806 : 1;
	8807 : 0;
	8808 : 0;
	8809 : 1;
	8810 : 1;
	8811 : 1;
	8812 : 1;
	8813 : 1;
	8814 : 1;
	8815 : 1;
	8816 : 1;
	8817 : 1;
	8818 : 1;
	8819 : 1;
	8820 : 1;
	8821 : 1;
	8822 : 0;
	8823 : 1;
	8824 : 1;
	8825 : 1;
	8826 : 1;
	8827 : 1;
	8828 : 1;
	8829 : 1;
	8830 : 1;
	8831 : 1;
	8832 : 1;
	8833 : 1;
	8834 : 1;
	8835 : 1;
	8836 : 1;
	8837 : 1;
	8838 : 1;
	8839 : 1;
	8840 : 1;
	8841 : 1;
	8842 : 1;
	8843 : 1;
	8844 : 1;
	8845 : 1;
	8846 : 1;
	8847 : 1;
	8848 : 1;
	8849 : 1;
	8850 : 1;
	8851 : 1;
	8852 : 1;
	8853 : 1;
	8854 : 1;
	8855 : 1;
	8856 : 1;
	8857 : 1;
	8858 : 1;
	8859 : 1;
	8860 : 1;
	8861 : 1;
	8862 : 1;
	8863 : 1;
	8864 : 1;
	8865 : 1;
	8866 : 1;
	8867 : 1;
	8868 : 1;
	8869 : 1;
	8870 : 1;
	8871 : 1;
	8872 : 1;
	8873 : 1;
	8874 : 1;
	8875 : 1;
	8876 : 1;
	8877 : 1;
	8878 : 1;
	8879 : 1;
	8880 : 1;
	8881 : 1;
	8882 : 1;
	8883 : 1;
	8884 : 1;
	8885 : 1;
	8886 : 1;
	8887 : 1;
	8888 : 1;
	8889 : 1;
	8890 : 1;
	8891 : 1;
	8892 : 1;
	8893 : 1;
	8894 : 1;
	8895 : 1;
	8896 : 1;
	8897 : 1;
	8898 : 1;
	8899 : 1;
	8900 : 1;
	8901 : 1;
	8902 : 1;
	8903 : 1;
	8904 : 1;
	8905 : 1;
	8906 : 1;
	8907 : 1;
	8908 : 1;
	8909 : 1;
	8910 : 1;
	8911 : 1;
	8912 : 1;
	8913 : 1;
	8914 : 1;
	8915 : 1;
	8916 : 1;
	8917 : 1;
	8918 : 1;
	8919 : 1;
	8920 : 1;
	8921 : 1;
	8922 : 1;
	8923 : 1;
	8924 : 1;
	8925 : 1;
	8926 : 1;
	8927 : 1;
	8928 : 1;
	8929 : 1;
	8930 : 1;
	8931 : 1;
	8932 : 1;
	8933 : 1;
	8934 : 1;
	8935 : 1;
	8936 : 0;
	8937 : 1;
	8938 : 1;
	8939 : 1;
	8940 : 0;
	8941 : 1;
	8942 : 0;
	8943 : 1;
	8944 : 1;
	8945 : 0;
	8946 : 0;
	8947 : 0;
	8948 : 0;
	8949 : 1;
	8950 : 1;
	8951 : 1;
	8952 : 0;
	8953 : 1;
	8954 : 1;
	8955 : 1;
	8956 : 0;
	8957 : 1;
	8958 : 1;
	8959 : 1;
	8960 : 0;
	8961 : 1;
	8962 : 0;
	8963 : 1;
	8964 : 1;
	8965 : 1;
	8966 : 0;
	8967 : 1;
	8968 : 0;
	8969 : 1;
	8970 : 1;
	8971 : 0;
	8972 : 0;
	8973 : 1;
	8974 : 0;
	8975 : 0;
	8976 : 0;
	8977 : 1;
	8978 : 1;
	8979 : 1;
	8980 : 1;
	8981 : 1;
	8982 : 0;
	8983 : 1;
	8984 : 1;
	8985 : 1;
	8986 : 1;
	8987 : 1;
	8988 : 0;
	8989 : 1;
	8990 : 0;
	8991 : 1;
	8992 : 1;
	8993 : 0;
	8994 : 0;
	8995 : 0;
	8996 : 1;
	8997 : 1;
	8998 : 1;
	8999 : 0;
	9000 : 0;
	9001 : 1;
	9002 : 0;
	9003 : 0;
	9004 : 1;
	9005 : 1;
	9006 : 1;
	9007 : 0;
	9008 : 0;
	9009 : 0;
	9010 : 0;
	9011 : 1;
	9012 : 1;
	9013 : 0;
	9014 : 0;
	9015 : 1;
	9016 : 1;
	9017 : 1;
	9018 : 0;
	9019 : 1;
	9020 : 1;
	9021 : 1;
	9022 : 0;
	9023 : 0;
	9024 : 1;
	9025 : 1;
	9026 : 1;
	9027 : 0;
	9028 : 0;
	9029 : 1;
	9030 : 0;
	9031 : 1;
	9032 : 1;
	9033 : 1;
	9034 : 0;
	9035 : 1;
	9036 : 0;
	9037 : 1;
	9038 : 1;
	9039 : 1;
	9040 : 0;
	9041 : 1;
	9042 : 1;
	9043 : 0;
	9044 : 1;
	9045 : 1;
	9046 : 1;
	9047 : 0;
	9048 : 0;
	9049 : 1;
	9050 : 1;
	9051 : 1;
	9052 : 1;
	9053 : 1;
	9054 : 1;
	9055 : 1;
	9056 : 1;
	9057 : 1;
	9058 : 1;
	9059 : 1;
	9060 : 1;
	9061 : 1;
	9062 : 0;
	9063 : 1;
	9064 : 1;
	9065 : 1;
	9066 : 1;
	9067 : 1;
	9068 : 1;
	9069 : 1;
	9070 : 1;
	9071 : 1;
	9072 : 1;
	9073 : 1;
	9074 : 1;
	9075 : 1;
	9076 : 1;
	9077 : 1;
	9078 : 1;
	9079 : 1;
	9080 : 1;
	9081 : 1;
	9082 : 1;
	9083 : 1;
	9084 : 1;
	9085 : 1;
	9086 : 1;
	9087 : 1;
	9088 : 1;
	9089 : 1;
	9090 : 1;
	9091 : 1;
	9092 : 1;
	9093 : 1;
	9094 : 1;
	9095 : 1;
	9096 : 1;
	9097 : 1;
	9098 : 1;
	9099 : 1;
	9100 : 1;
	9101 : 1;
	9102 : 1;
	9103 : 1;
	9104 : 1;
	9105 : 1;
	9106 : 1;
	9107 : 1;
	9108 : 1;
	9109 : 1;
	9110 : 1;
	9111 : 1;
	9112 : 1;
	9113 : 1;
	9114 : 1;
	9115 : 1;
	9116 : 1;
	9117 : 1;
	9118 : 1;
	9119 : 1;
	9120 : 1;
	9121 : 1;
	9122 : 1;
	9123 : 1;
	9124 : 1;
	9125 : 1;
	9126 : 1;
	9127 : 1;
	9128 : 1;
	9129 : 1;
	9130 : 1;
	9131 : 1;
	9132 : 1;
	9133 : 1;
	9134 : 1;
	9135 : 1;
	9136 : 1;
	9137 : 1;
	9138 : 1;
	9139 : 1;
	9140 : 1;
	9141 : 1;
	9142 : 1;
	9143 : 1;
	9144 : 1;
	9145 : 1;
	9146 : 1;
	9147 : 1;
	9148 : 1;
	9149 : 1;
	9150 : 1;
	9151 : 1;
	9152 : 1;
	9153 : 1;
	9154 : 1;
	9155 : 1;
	9156 : 1;
	9157 : 1;
	9158 : 1;
	9159 : 1;
	9160 : 1;
	9161 : 1;
	9162 : 1;
	9163 : 1;
	9164 : 1;
	9165 : 1;
	9166 : 1;
	9167 : 1;
	9168 : 1;
	9169 : 1;
	9170 : 1;
	9171 : 1;
	9172 : 1;
	9173 : 1;
	9174 : 1;
	9175 : 1;
	9176 : 0;
	9177 : 1;
	9178 : 1;
	9179 : 1;
	9180 : 0;
	9181 : 1;
	9182 : 0;
	9183 : 1;
	9184 : 1;
	9185 : 0;
	9186 : 0;
	9187 : 0;
	9188 : 0;
	9189 : 1;
	9190 : 1;
	9191 : 1;
	9192 : 0;
	9193 : 1;
	9194 : 1;
	9195 : 1;
	9196 : 0;
	9197 : 1;
	9198 : 1;
	9199 : 1;
	9200 : 0;
	9201 : 1;
	9202 : 0;
	9203 : 1;
	9204 : 1;
	9205 : 1;
	9206 : 0;
	9207 : 1;
	9208 : 0;
	9209 : 1;
	9210 : 1;
	9211 : 0;
	9212 : 0;
	9213 : 1;
	9214 : 0;
	9215 : 0;
	9216 : 1;
	9217 : 1;
	9218 : 1;
	9219 : 1;
	9220 : 1;
	9221 : 1;
	9222 : 0;
	9223 : 1;
	9224 : 1;
	9225 : 1;
	9226 : 1;
	9227 : 1;
	9228 : 0;
	9229 : 1;
	9230 : 0;
	9231 : 1;
	9232 : 1;
	9233 : 0;
	9234 : 0;
	9235 : 0;
	9236 : 1;
	9237 : 1;
	9238 : 1;
	9239 : 0;
	9240 : 0;
	9241 : 1;
	9242 : 0;
	9243 : 0;
	9244 : 1;
	9245 : 1;
	9246 : 1;
	9247 : 0;
	9248 : 1;
	9249 : 1;
	9250 : 1;
	9251 : 1;
	9252 : 1;
	9253 : 0;
	9254 : 1;
	9255 : 1;
	9256 : 1;
	9257 : 1;
	9258 : 0;
	9259 : 1;
	9260 : 1;
	9261 : 1;
	9262 : 0;
	9263 : 0;
	9264 : 1;
	9265 : 1;
	9266 : 1;
	9267 : 0;
	9268 : 0;
	9269 : 1;
	9270 : 0;
	9271 : 0;
	9272 : 0;
	9273 : 0;
	9274 : 0;
	9275 : 1;
	9276 : 0;
	9277 : 1;
	9278 : 1;
	9279 : 1;
	9280 : 1;
	9281 : 1;
	9282 : 1;
	9283 : 0;
	9284 : 1;
	9285 : 1;
	9286 : 1;
	9287 : 1;
	9288 : 1;
	9289 : 1;
	9290 : 1;
	9291 : 1;
	9292 : 1;
	9293 : 1;
	9294 : 1;
	9295 : 1;
	9296 : 1;
	9297 : 1;
	9298 : 0;
	9299 : 0;
	9300 : 1;
	9301 : 1;
	9302 : 0;
	9303 : 1;
	9304 : 1;
	9305 : 1;
	9306 : 1;
	9307 : 1;
	9308 : 1;
	9309 : 1;
	9310 : 1;
	9311 : 1;
	9312 : 1;
	9313 : 1;
	9314 : 1;
	9315 : 1;
	9316 : 1;
	9317 : 1;
	9318 : 1;
	9319 : 1;
	9320 : 1;
	9321 : 1;
	9322 : 1;
	9323 : 1;
	9324 : 1;
	9325 : 1;
	9326 : 1;
	9327 : 1;
	9328 : 1;
	9329 : 1;
	9330 : 1;
	9331 : 1;
	9332 : 1;
	9333 : 1;
	9334 : 1;
	9335 : 1;
	9336 : 1;
	9337 : 1;
	9338 : 1;
	9339 : 1;
	9340 : 1;
	9341 : 1;
	9342 : 1;
	9343 : 1;
	9344 : 1;
	9345 : 1;
	9346 : 1;
	9347 : 1;
	9348 : 1;
	9349 : 1;
	9350 : 1;
	9351 : 1;
	9352 : 1;
	9353 : 1;
	9354 : 1;
	9355 : 1;
	9356 : 1;
	9357 : 1;
	9358 : 1;
	9359 : 1;
	9360 : 1;
	9361 : 1;
	9362 : 1;
	9363 : 1;
	9364 : 1;
	9365 : 1;
	9366 : 1;
	9367 : 1;
	9368 : 1;
	9369 : 1;
	9370 : 1;
	9371 : 1;
	9372 : 1;
	9373 : 1;
	9374 : 1;
	9375 : 1;
	9376 : 1;
	9377 : 1;
	9378 : 1;
	9379 : 1;
	9380 : 1;
	9381 : 1;
	9382 : 1;
	9383 : 1;
	9384 : 1;
	9385 : 1;
	9386 : 1;
	9387 : 1;
	9388 : 1;
	9389 : 1;
	9390 : 1;
	9391 : 1;
	9392 : 1;
	9393 : 1;
	9394 : 1;
	9395 : 1;
	9396 : 1;
	9397 : 1;
	9398 : 1;
	9399 : 1;
	9400 : 1;
	9401 : 1;
	9402 : 1;
	9403 : 1;
	9404 : 1;
	9405 : 1;
	9406 : 1;
	9407 : 1;
	9408 : 1;
	9409 : 1;
	9410 : 1;
	9411 : 1;
	9412 : 1;
	9413 : 1;
	9414 : 1;
	9415 : 1;
	9416 : 0;
	9417 : 1;
	9418 : 1;
	9419 : 0;
	9420 : 0;
	9421 : 1;
	9422 : 0;
	9423 : 1;
	9424 : 1;
	9425 : 0;
	9426 : 0;
	9427 : 0;
	9428 : 0;
	9429 : 1;
	9430 : 1;
	9431 : 1;
	9432 : 0;
	9433 : 1;
	9434 : 1;
	9435 : 1;
	9436 : 0;
	9437 : 1;
	9438 : 1;
	9439 : 1;
	9440 : 0;
	9441 : 1;
	9442 : 0;
	9443 : 1;
	9444 : 1;
	9445 : 1;
	9446 : 0;
	9447 : 1;
	9448 : 0;
	9449 : 1;
	9450 : 1;
	9451 : 0;
	9452 : 0;
	9453 : 1;
	9454 : 0;
	9455 : 0;
	9456 : 1;
	9457 : 1;
	9458 : 1;
	9459 : 1;
	9460 : 1;
	9461 : 1;
	9462 : 0;
	9463 : 1;
	9464 : 1;
	9465 : 1;
	9466 : 1;
	9467 : 1;
	9468 : 0;
	9469 : 1;
	9470 : 0;
	9471 : 1;
	9472 : 1;
	9473 : 0;
	9474 : 0;
	9475 : 0;
	9476 : 1;
	9477 : 1;
	9478 : 0;
	9479 : 0;
	9480 : 0;
	9481 : 1;
	9482 : 0;
	9483 : 0;
	9484 : 1;
	9485 : 1;
	9486 : 1;
	9487 : 0;
	9488 : 1;
	9489 : 1;
	9490 : 1;
	9491 : 1;
	9492 : 1;
	9493 : 0;
	9494 : 1;
	9495 : 1;
	9496 : 1;
	9497 : 1;
	9498 : 0;
	9499 : 1;
	9500 : 1;
	9501 : 1;
	9502 : 0;
	9503 : 0;
	9504 : 1;
	9505 : 1;
	9506 : 1;
	9507 : 0;
	9508 : 0;
	9509 : 1;
	9510 : 0;
	9511 : 1;
	9512 : 1;
	9513 : 1;
	9514 : 1;
	9515 : 1;
	9516 : 0;
	9517 : 1;
	9518 : 1;
	9519 : 1;
	9520 : 0;
	9521 : 1;
	9522 : 1;
	9523 : 0;
	9524 : 1;
	9525 : 1;
	9526 : 1;
	9527 : 0;
	9528 : 0;
	9529 : 1;
	9530 : 1;
	9531 : 1;
	9532 : 1;
	9533 : 1;
	9534 : 1;
	9535 : 1;
	9536 : 1;
	9537 : 1;
	9538 : 0;
	9539 : 0;
	9540 : 1;
	9541 : 1;
	9542 : 0;
	9543 : 1;
	9544 : 1;
	9545 : 1;
	9546 : 1;
	9547 : 1;
	9548 : 1;
	9549 : 1;
	9550 : 1;
	9551 : 1;
	9552 : 1;
	9553 : 1;
	9554 : 1;
	9555 : 1;
	9556 : 1;
	9557 : 1;
	9558 : 1;
	9559 : 1;
	9560 : 1;
	9561 : 1;
	9562 : 1;
	9563 : 1;
	9564 : 1;
	9565 : 1;
	9566 : 1;
	9567 : 1;
	9568 : 1;
	9569 : 1;
	9570 : 1;
	9571 : 1;
	9572 : 1;
	9573 : 1;
	9574 : 1;
	9575 : 1;
	9576 : 1;
	9577 : 1;
	9578 : 1;
	9579 : 1;
	9580 : 1;
	9581 : 1;
	9582 : 1;
	9583 : 1;
	9584 : 1;
	9585 : 1;
	9586 : 1;
	9587 : 1;
	9588 : 1;
	9589 : 1;
	9590 : 1;
	9591 : 1;
	9592 : 1;
	9593 : 1;
	9594 : 1;
	9595 : 1;
	9596 : 1;
	9597 : 1;
	9598 : 1;
	9599 : 1;
	9600 : 1;
	9601 : 1;
	9602 : 1;
	9603 : 1;
	9604 : 1;
	9605 : 1;
	9606 : 1;
	9607 : 1;
	9608 : 1;
	9609 : 1;
	9610 : 1;
	9611 : 1;
	9612 : 1;
	9613 : 1;
	9614 : 1;
	9615 : 1;
	9616 : 1;
	9617 : 1;
	9618 : 1;
	9619 : 1;
	9620 : 1;
	9621 : 1;
	9622 : 1;
	9623 : 1;
	9624 : 1;
	9625 : 1;
	9626 : 1;
	9627 : 1;
	9628 : 1;
	9629 : 1;
	9630 : 1;
	9631 : 1;
	9632 : 1;
	9633 : 1;
	9634 : 1;
	9635 : 1;
	9636 : 1;
	9637 : 1;
	9638 : 1;
	9639 : 1;
	9640 : 1;
	9641 : 1;
	9642 : 1;
	9643 : 1;
	9644 : 1;
	9645 : 1;
	9646 : 1;
	9647 : 1;
	9648 : 1;
	9649 : 1;
	9650 : 1;
	9651 : 1;
	9652 : 1;
	9653 : 1;
	9654 : 1;
	9655 : 1;
	9656 : 1;
	9657 : 0;
	9658 : 0;
	9659 : 1;
	9660 : 0;
	9661 : 1;
	9662 : 0;
	9663 : 1;
	9664 : 1;
	9665 : 0;
	9666 : 0;
	9667 : 1;
	9668 : 0;
	9669 : 0;
	9670 : 0;
	9671 : 0;
	9672 : 0;
	9673 : 1;
	9674 : 1;
	9675 : 1;
	9676 : 1;
	9677 : 0;
	9678 : 0;
	9679 : 0;
	9680 : 0;
	9681 : 1;
	9682 : 1;
	9683 : 0;
	9684 : 0;
	9685 : 0;
	9686 : 1;
	9687 : 1;
	9688 : 1;
	9689 : 0;
	9690 : 0;
	9691 : 0;
	9692 : 0;
	9693 : 0;
	9694 : 0;
	9695 : 0;
	9696 : 1;
	9697 : 1;
	9698 : 1;
	9699 : 1;
	9700 : 1;
	9701 : 1;
	9702 : 0;
	9703 : 1;
	9704 : 1;
	9705 : 1;
	9706 : 1;
	9707 : 1;
	9708 : 0;
	9709 : 1;
	9710 : 0;
	9711 : 1;
	9712 : 1;
	9713 : 0;
	9714 : 0;
	9715 : 1;
	9716 : 0;
	9717 : 0;
	9718 : 0;
	9719 : 0;
	9720 : 0;
	9721 : 1;
	9722 : 0;
	9723 : 0;
	9724 : 1;
	9725 : 1;
	9726 : 1;
	9727 : 0;
	9728 : 1;
	9729 : 1;
	9730 : 1;
	9731 : 1;
	9732 : 1;
	9733 : 0;
	9734 : 1;
	9735 : 1;
	9736 : 1;
	9737 : 1;
	9738 : 1;
	9739 : 0;
	9740 : 0;
	9741 : 0;
	9742 : 0;
	9743 : 1;
	9744 : 0;
	9745 : 0;
	9746 : 1;
	9747 : 0;
	9748 : 0;
	9749 : 1;
	9750 : 1;
	9751 : 0;
	9752 : 0;
	9753 : 0;
	9754 : 0;
	9755 : 1;
	9756 : 1;
	9757 : 0;
	9758 : 0;
	9759 : 0;
	9760 : 1;
	9761 : 1;
	9762 : 1;
	9763 : 0;
	9764 : 0;
	9765 : 0;
	9766 : 0;
	9767 : 0;
	9768 : 0;
	9769 : 1;
	9770 : 1;
	9771 : 1;
	9772 : 1;
	9773 : 1;
	9774 : 1;
	9775 : 1;
	9776 : 1;
	9777 : 1;
	9778 : 1;
	9779 : 0;
	9780 : 1;
	9781 : 0;
	9782 : 1;
	9783 : 1;
	9784 : 1;
	9785 : 1;
	9786 : 1;
	9787 : 1;
	9788 : 1;
	9789 : 1;
	9790 : 1;
	9791 : 1;
	9792 : 1;
	9793 : 1;
	9794 : 1;
	9795 : 1;
	9796 : 1;
	9797 : 1;
	9798 : 1;
	9799 : 1;
	9800 : 1;
	9801 : 1;
	9802 : 1;
	9803 : 1;
	9804 : 1;
	9805 : 1;
	9806 : 1;
	9807 : 1;
	9808 : 1;
	9809 : 1;
	9810 : 1;
	9811 : 1;
	9812 : 1;
	9813 : 1;
	9814 : 1;
	9815 : 1;
	9816 : 1;
	9817 : 1;
	9818 : 1;
	9819 : 1;
	9820 : 1;
	9821 : 1;
	9822 : 1;
	9823 : 1;
	9824 : 1;
	9825 : 1;
	9826 : 1;
	9827 : 1;
	9828 : 1;
	9829 : 1;
	9830 : 1;
	9831 : 1;
	9832 : 1;
	9833 : 1;
	9834 : 1;
	9835 : 1;
	9836 : 1;
	9837 : 1;
	9838 : 1;
	9839 : 1;
	9840 : 1;
	9841 : 1;
	9842 : 1;
	9843 : 1;
	9844 : 1;
	9845 : 1;
	9846 : 1;
	9847 : 1;
	9848 : 1;
	9849 : 1;
	9850 : 1;
	9851 : 1;
	9852 : 1;
	9853 : 1;
	9854 : 1;
	9855 : 1;
	9856 : 1;
	9857 : 1;
	9858 : 1;
	9859 : 1;
	9860 : 1;
	9861 : 1;
	9862 : 1;
	9863 : 1;
	9864 : 1;
	9865 : 1;
	9866 : 1;
	9867 : 1;
	9868 : 1;
	9869 : 1;
	9870 : 1;
	9871 : 1;
	9872 : 1;
	9873 : 1;
	9874 : 1;
	9875 : 1;
	9876 : 1;
	9877 : 1;
	9878 : 1;
	9879 : 1;
	9880 : 1;
	9881 : 1;
	9882 : 1;
	9883 : 1;
	9884 : 1;
	9885 : 1;
	9886 : 1;
	9887 : 1;
	9888 : 1;
	9889 : 1;
	9890 : 1;
	9891 : 1;
	9892 : 1;
	9893 : 1;
	9894 : 1;
	9895 : 1;
	9896 : 1;
	9897 : 1;
	9898 : 1;
	9899 : 1;
	9900 : 1;
	9901 : 1;
	9902 : 1;
	9903 : 1;
	9904 : 1;
	9905 : 1;
	9906 : 1;
	9907 : 1;
	9908 : 1;
	9909 : 1;
	9910 : 1;
	9911 : 1;
	9912 : 1;
	9913 : 1;
	9914 : 1;
	9915 : 1;
	9916 : 1;
	9917 : 1;
	9918 : 1;
	9919 : 1;
	9920 : 0;
	9921 : 1;
	9922 : 1;
	9923 : 1;
	9924 : 1;
	9925 : 1;
	9926 : 1;
	9927 : 1;
	9928 : 1;
	9929 : 1;
	9930 : 1;
	9931 : 1;
	9932 : 1;
	9933 : 1;
	9934 : 1;
	9935 : 1;
	9936 : 1;
	9937 : 1;
	9938 : 1;
	9939 : 1;
	9940 : 1;
	9941 : 1;
	9942 : 1;
	9943 : 1;
	9944 : 1;
	9945 : 1;
	9946 : 1;
	9947 : 1;
	9948 : 1;
	9949 : 1;
	9950 : 1;
	9951 : 1;
	9952 : 1;
	9953 : 1;
	9954 : 1;
	9955 : 1;
	9956 : 1;
	9957 : 1;
	9958 : 1;
	9959 : 1;
	9960 : 1;
	9961 : 1;
	9962 : 1;
	9963 : 1;
	9964 : 1;
	9965 : 1;
	9966 : 1;
	9967 : 1;
	9968 : 1;
	9969 : 1;
	9970 : 1;
	9971 : 1;
	9972 : 1;
	9973 : 1;
	9974 : 1;
	9975 : 1;
	9976 : 1;
	9977 : 1;
	9978 : 1;
	9979 : 1;
	9980 : 1;
	9981 : 1;
	9982 : 1;
	9983 : 1;
	9984 : 0;
	9985 : 0;
	9986 : 1;
	9987 : 0;
	9988 : 0;
	9989 : 1;
	9990 : 1;
	9991 : 1;
	9992 : 1;
	9993 : 1;
	9994 : 1;
	9995 : 1;
	9996 : 1;
	9997 : 1;
	9998 : 1;
	9999 : 1;
	10000 : 1;
	10001 : 1;
	10002 : 1;
	10003 : 1;
	10004 : 1;
	10005 : 1;
	10006 : 1;
	10007 : 1;
	10008 : 1;
	10009 : 1;
	10010 : 1;
	10011 : 1;
	10012 : 1;
	10013 : 1;
	10014 : 1;
	10015 : 1;
	10016 : 1;
	10017 : 1;
	10018 : 0;
	10019 : 1;
	10020 : 1;
	10021 : 1;
	10022 : 1;
	10023 : 1;
	10024 : 1;
	10025 : 1;
	10026 : 1;
	10027 : 1;
	10028 : 1;
	10029 : 1;
	10030 : 1;
	10031 : 1;
	10032 : 1;
	10033 : 1;
	10034 : 1;
	10035 : 1;
	10036 : 1;
	10037 : 1;
	10038 : 1;
	10039 : 1;
	10040 : 1;
	10041 : 1;
	10042 : 1;
	10043 : 1;
	10044 : 1;
	10045 : 1;
	10046 : 1;
	10047 : 1;
	10048 : 1;
	10049 : 1;
	10050 : 1;
	10051 : 1;
	10052 : 1;
	10053 : 1;
	10054 : 1;
	10055 : 1;
	10056 : 1;
	10057 : 1;
	10058 : 1;
	10059 : 1;
	10060 : 1;
	10061 : 1;
	10062 : 1;
	10063 : 1;
	10064 : 1;
	10065 : 1;
	10066 : 1;
	10067 : 1;
	10068 : 1;
	10069 : 1;
	10070 : 1;
	10071 : 1;
	10072 : 1;
	10073 : 1;
	10074 : 1;
	10075 : 1;
	10076 : 1;
	10077 : 1;
	10078 : 1;
	10079 : 1;
	10080 : 1;
	10081 : 1;
	10082 : 1;
	10083 : 1;
	10084 : 1;
	10085 : 1;
	10086 : 1;
	10087 : 1;
	10088 : 1;
	10089 : 1;
	10090 : 1;
	10091 : 1;
	10092 : 1;
	10093 : 1;
	10094 : 1;
	10095 : 1;
	10096 : 1;
	10097 : 1;
	10098 : 1;
	10099 : 1;
	10100 : 1;
	10101 : 1;
	10102 : 1;
	10103 : 1;
	10104 : 1;
	10105 : 1;
	10106 : 1;
	10107 : 1;
	10108 : 1;
	10109 : 1;
	10110 : 1;
	10111 : 1;
	10112 : 1;
	10113 : 1;
	10114 : 1;
	10115 : 1;
	10116 : 1;
	10117 : 1;
	10118 : 1;
	10119 : 1;
	10120 : 1;
	10121 : 1;
	10122 : 1;
	10123 : 1;
	10124 : 1;
	10125 : 1;
	10126 : 1;
	10127 : 1;
	10128 : 1;
	10129 : 1;
	10130 : 1;
	10131 : 1;
	10132 : 1;
	10133 : 1;
	10134 : 1;
	10135 : 1;
	10136 : 1;
	10137 : 1;
	10138 : 1;
	10139 : 1;
	10140 : 1;
	10141 : 1;
	10142 : 1;
	10143 : 1;
	10144 : 1;
	10145 : 1;
	10146 : 1;
	10147 : 1;
	10148 : 1;
	10149 : 1;
	10150 : 1;
	10151 : 1;
	10152 : 1;
	10153 : 1;
	10154 : 1;
	10155 : 1;
	10156 : 0;
	10157 : 0;
	10158 : 0;
	10159 : 0;
	10160 : 1;
	10161 : 1;
	10162 : 1;
	10163 : 1;
	10164 : 1;
	10165 : 1;
	10166 : 1;
	10167 : 1;
	10168 : 1;
	10169 : 1;
	10170 : 1;
	10171 : 1;
	10172 : 1;
	10173 : 1;
	10174 : 1;
	10175 : 1;
	10176 : 1;
	10177 : 1;
	10178 : 1;
	10179 : 1;
	10180 : 1;
	10181 : 1;
	10182 : 1;
	10183 : 1;
	10184 : 1;
	10185 : 1;
	10186 : 1;
	10187 : 1;
	10188 : 1;
	10189 : 1;
	10190 : 1;
	10191 : 1;
	10192 : 1;
	10193 : 1;
	10194 : 1;
	10195 : 1;
	10196 : 1;
	10197 : 1;
	10198 : 1;
	10199 : 1;
	10200 : 1;
	10201 : 1;
	10202 : 1;
	10203 : 1;
	10204 : 1;
	10205 : 1;
	10206 : 1;
	10207 : 1;
	10208 : 1;
	10209 : 1;
	10210 : 1;
	10211 : 1;
	10212 : 1;
	10213 : 1;
	10214 : 1;
	10215 : 1;
	10216 : 1;
	10217 : 1;
	10218 : 1;
	10219 : 1;
	10220 : 1;
	10221 : 1;
	10222 : 1;
	10223 : 1;
	10224 : 1;
	10225 : 0;
	10226 : 0;
	10227 : 0;
	10228 : 1;
	10229 : 1;
	10230 : 1;
	10231 : 1;
	10232 : 1;
	10233 : 1;
	10234 : 1;
	10235 : 1;
	10236 : 1;
	10237 : 1;
	10238 : 1;
	10239 : 1;
	10240 : 1;
	10241 : 1;
	10242 : 1;
	10243 : 1;
	10244 : 1;
	10245 : 1;
	10246 : 1;
	10247 : 1;
	10248 : 1;
	10249 : 1;
	10250 : 1;
	10251 : 1;
	10252 : 1;
	10253 : 1;
	10254 : 1;
	10255 : 1;
	10256 : 1;
	10257 : 1;
	10258 : 1;
	10259 : 1;
	10260 : 1;
	10261 : 1;
	10262 : 1;
	10263 : 1;
	10264 : 1;
	10265 : 1;
	10266 : 1;
	10267 : 1;
	10268 : 1;
	10269 : 1;
	10270 : 1;
	10271 : 1;
	10272 : 1;
	10273 : 1;
	10274 : 1;
	10275 : 1;
	10276 : 1;
	10277 : 1;
	10278 : 1;
	10279 : 1;
	10280 : 1;
	10281 : 1;
	10282 : 1;
	10283 : 1;
	10284 : 1;
	10285 : 1;
	10286 : 1;
	10287 : 1;
	10288 : 1;
	10289 : 1;
	10290 : 1;
	10291 : 1;
	10292 : 1;
	10293 : 1;
	10294 : 1;
	10295 : 1;
	10296 : 1;
	10297 : 1;
	10298 : 1;
	10299 : 1;
	10300 : 1;
	10301 : 1;
	10302 : 1;
	10303 : 1;
	10304 : 1;
	10305 : 1;
	10306 : 1;
	10307 : 1;
	10308 : 1;
	10309 : 1;
	10310 : 1;
	10311 : 1;
	10312 : 1;
	10313 : 1;
	10314 : 1;
	10315 : 1;
	10316 : 1;
	10317 : 1;
	10318 : 1;
	10319 : 1;
	10320 : 1;
	10321 : 1;
	10322 : 1;
	10323 : 1;
	10324 : 1;
	10325 : 1;
	10326 : 1;
	10327 : 1;
	10328 : 1;
	10329 : 1;
	10330 : 1;
	10331 : 1;
	10332 : 1;
	10333 : 1;
	10334 : 1;
	10335 : 1;
	10336 : 1;
	10337 : 1;
	10338 : 1;
	10339 : 1;
	10340 : 1;
	10341 : 1;
	10342 : 1;
	10343 : 1;
	10344 : 1;
	10345 : 1;
	10346 : 1;
	10347 : 1;
	10348 : 1;
	10349 : 1;
	10350 : 1;
	10351 : 1;
	10352 : 1;
	10353 : 1;
	10354 : 1;
	10355 : 1;
	10356 : 1;
	10357 : 1;
	10358 : 1;
	10359 : 1;
	10360 : 1;
	10361 : 1;
	10362 : 1;
	10363 : 1;
	10364 : 1;
	10365 : 1;
	10366 : 1;
	10367 : 1;
	10368 : 1;
	10369 : 1;
	10370 : 1;
	10371 : 1;
	10372 : 1;
	10373 : 1;
	10374 : 1;
	10375 : 1;
	10376 : 1;
	10377 : 1;
	10378 : 1;
	10379 : 1;
	10380 : 1;
	10381 : 1;
	10382 : 1;
	10383 : 1;
	10384 : 1;
	10385 : 1;
	10386 : 1;
	10387 : 1;
	10388 : 1;
	10389 : 1;
	10390 : 1;
	10391 : 1;
	10392 : 1;
	10393 : 1;
	10394 : 1;
	10395 : 1;
	10396 : 1;
	10397 : 1;
	10398 : 1;
	10399 : 1;
	10400 : 1;
	10401 : 1;
	10402 : 1;
	10403 : 1;
	10404 : 1;
	10405 : 1;
	10406 : 1;
	10407 : 1;
	10408 : 1;
	10409 : 1;
	10410 : 1;
	10411 : 1;
	10412 : 1;
	10413 : 1;
	10414 : 1;
	10415 : 1;
	10416 : 1;
	10417 : 1;
	10418 : 1;
	10419 : 1;
	10420 : 1;
	10421 : 1;
	10422 : 1;
	10423 : 1;
	10424 : 1;
	10425 : 1;
	10426 : 1;
	10427 : 1;
	10428 : 1;
	10429 : 1;
	10430 : 1;
	10431 : 1;
	10432 : 1;
	10433 : 1;
	10434 : 1;
	10435 : 1;
	10436 : 1;
	10437 : 1;
	10438 : 1;
	10439 : 1;
	10440 : 1;
	10441 : 1;
	10442 : 1;
	10443 : 1;
	10444 : 1;
	10445 : 1;
	10446 : 1;
	10447 : 1;
	10448 : 1;
	10449 : 1;
	10450 : 1;
	10451 : 1;
	10452 : 1;
	10453 : 1;
	10454 : 1;
	10455 : 1;
	10456 : 1;
	10457 : 1;
	10458 : 1;
	10459 : 1;
	10460 : 1;
	10461 : 1;
	10462 : 1;
	10463 : 1;
	10464 : 1;
	10465 : 1;
	10466 : 1;
	10467 : 1;
	10468 : 1;
	10469 : 1;
	10470 : 1;
	10471 : 1;
	10472 : 1;
	10473 : 1;
	10474 : 1;
	10475 : 1;
	10476 : 1;
	10477 : 1;
	10478 : 1;
	10479 : 1;
	10480 : 1;
	10481 : 1;
	10482 : 1;
	10483 : 1;
	10484 : 1;
	10485 : 1;
	10486 : 1;
	10487 : 1;
	10488 : 1;
	10489 : 1;
	10490 : 1;
	10491 : 1;
	10492 : 1;
	10493 : 1;
	10494 : 1;
	10495 : 1;
	10496 : 1;
	10497 : 1;
	10498 : 1;
	10499 : 1;
	10500 : 1;
	10501 : 1;
	10502 : 1;
	10503 : 1;
	10504 : 1;
	10505 : 1;
	10506 : 1;
	10507 : 1;
	10508 : 1;
	10509 : 1;
	10510 : 1;
	10511 : 1;
	10512 : 1;
	10513 : 1;
	10514 : 1;
	10515 : 1;
	10516 : 1;
	10517 : 1;
	10518 : 1;
	10519 : 1;
	10520 : 1;
	10521 : 1;
	10522 : 1;
	10523 : 1;
	10524 : 1;
	10525 : 1;
	10526 : 1;
	10527 : 1;
	10528 : 1;
	10529 : 1;
	10530 : 1;
	10531 : 1;
	10532 : 1;
	10533 : 1;
	10534 : 1;
	10535 : 1;
	10536 : 1;
	10537 : 1;
	10538 : 1;
	10539 : 1;
	10540 : 1;
	10541 : 1;
	10542 : 1;
	10543 : 1;
	10544 : 1;
	10545 : 1;
	10546 : 1;
	10547 : 1;
	10548 : 1;
	10549 : 1;
	10550 : 1;
	10551 : 1;
	10552 : 1;
	10553 : 1;
	10554 : 1;
	10555 : 1;
	10556 : 1;
	10557 : 1;
	10558 : 1;
	10559 : 1;
	10560 : 1;
	10561 : 1;
	10562 : 1;
	10563 : 1;
	10564 : 1;
	10565 : 1;
	10566 : 1;
	10567 : 1;
	10568 : 1;
	10569 : 1;
	10570 : 1;
	10571 : 1;
	10572 : 1;
	10573 : 1;
	10574 : 1;
	10575 : 1;
	10576 : 1;
	10577 : 1;
	10578 : 1;
	10579 : 1;
	10580 : 1;
	10581 : 1;
	10582 : 1;
	10583 : 1;
	10584 : 1;
	10585 : 1;
	10586 : 1;
	10587 : 1;
	10588 : 1;
	10589 : 1;
	10590 : 1;
	10591 : 1;
	10592 : 1;
	10593 : 1;
	10594 : 1;
	10595 : 1;
	10596 : 1;
	10597 : 1;
	10598 : 1;
	10599 : 1;
	10600 : 1;
	10601 : 1;
	10602 : 1;
	10603 : 1;
	10604 : 1;
	10605 : 1;
	10606 : 1;
	10607 : 1;
	10608 : 1;
	10609 : 1;
	10610 : 1;
	10611 : 1;
	10612 : 1;
	10613 : 1;
	10614 : 1;
	10615 : 1;
	10616 : 1;
	10617 : 1;
	10618 : 1;
	10619 : 1;
	10620 : 1;
	10621 : 1;
	10622 : 1;
	10623 : 1;
	10624 : 1;
	10625 : 1;
	10626 : 1;
	10627 : 1;
	10628 : 1;
	10629 : 1;
	10630 : 1;
	10631 : 1;
	10632 : 1;
	10633 : 1;
	10634 : 1;
	10635 : 1;
	10636 : 1;
	10637 : 1;
	10638 : 1;
	10639 : 1;
	10640 : 1;
	10641 : 1;
	10642 : 1;
	10643 : 1;
	10644 : 1;
	10645 : 1;
	10646 : 1;
	10647 : 1;
	10648 : 1;
	10649 : 1;
	10650 : 1;
	10651 : 1;
	10652 : 1;
	10653 : 1;
	10654 : 1;
	10655 : 1;
	10656 : 1;
	10657 : 1;
	10658 : 1;
	10659 : 1;
	10660 : 1;
	10661 : 1;
	10662 : 1;
	10663 : 1;
	10664 : 1;
	10665 : 1;
	10666 : 1;
	10667 : 1;
	10668 : 1;
	10669 : 1;
	10670 : 1;
	10671 : 1;
	10672 : 1;
	10673 : 1;
	10674 : 1;
	10675 : 1;
	10676 : 1;
	10677 : 1;
	10678 : 1;
	10679 : 1;
	10680 : 1;
	10681 : 1;
	10682 : 1;
	10683 : 1;
	10684 : 1;
	10685 : 1;
	10686 : 1;
	10687 : 1;
	10688 : 1;
	10689 : 1;
	10690 : 1;
	10691 : 1;
	10692 : 1;
	10693 : 1;
	10694 : 1;
	10695 : 1;
	10696 : 1;
	10697 : 1;
	10698 : 1;
	10699 : 1;
	10700 : 1;
	10701 : 1;
	10702 : 1;
	10703 : 1;
	10704 : 1;
	10705 : 1;
	10706 : 1;
	10707 : 1;
	10708 : 1;
	10709 : 1;
	10710 : 1;
	10711 : 1;
	10712 : 1;
	10713 : 1;
	10714 : 1;
	10715 : 1;
	10716 : 1;
	10717 : 1;
	10718 : 1;
	10719 : 1;
	10720 : 1;
	10721 : 1;
	10722 : 1;
	10723 : 1;
	10724 : 1;
	10725 : 1;
	10726 : 1;
	10727 : 1;
	10728 : 1;
	10729 : 1;
	10730 : 1;
	10731 : 1;
	10732 : 1;
	10733 : 1;
	10734 : 1;
	10735 : 1;
	10736 : 1;
	10737 : 1;
	10738 : 1;
	10739 : 1;
	10740 : 1;
	10741 : 1;
	10742 : 1;
	10743 : 1;
	10744 : 1;
	10745 : 1;
	10746 : 1;
	10747 : 1;
	10748 : 1;
	10749 : 1;
	10750 : 1;
	10751 : 1;
	10752 : 1;
	10753 : 1;
	10754 : 1;
	10755 : 1;
	10756 : 1;
	10757 : 1;
	10758 : 1;
	10759 : 1;
	10760 : 1;
	10761 : 1;
	10762 : 1;
	10763 : 1;
	10764 : 1;
	10765 : 1;
	10766 : 1;
	10767 : 1;
	10768 : 1;
	10769 : 1;
	10770 : 1;
	10771 : 1;
	10772 : 1;
	10773 : 1;
	10774 : 1;
	10775 : 1;
	10776 : 1;
	10777 : 1;
	10778 : 1;
	10779 : 1;
	10780 : 1;
	10781 : 1;
	10782 : 1;
	10783 : 1;
	10784 : 1;
	10785 : 1;
	10786 : 1;
	10787 : 1;
	10788 : 1;
	10789 : 1;
	10790 : 1;
	10791 : 1;
	10792 : 1;
	10793 : 1;
	10794 : 1;
	10795 : 1;
	10796 : 1;
	10797 : 1;
	10798 : 1;
	10799 : 1;
	10800 : 1;
	10801 : 1;
	10802 : 1;
	10803 : 1;
	10804 : 1;
	10805 : 1;
	10806 : 1;
	10807 : 1;
	10808 : 1;
	10809 : 1;
	10810 : 1;
	10811 : 1;
	10812 : 1;
	10813 : 1;
	10814 : 1;
	10815 : 1;
	10816 : 1;
	10817 : 1;
	10818 : 1;
	10819 : 1;
	10820 : 1;
	10821 : 1;
	10822 : 1;
	10823 : 1;
	10824 : 1;
	10825 : 1;
	10826 : 1;
	10827 : 1;
	10828 : 1;
	10829 : 1;
	10830 : 1;
	10831 : 1;
	10832 : 1;
	10833 : 1;
	10834 : 1;
	10835 : 1;
	10836 : 1;
	10837 : 1;
	10838 : 1;
	10839 : 1;
	10840 : 1;
	10841 : 1;
	10842 : 1;
	10843 : 1;
	10844 : 1;
	10845 : 1;
	10846 : 1;
	10847 : 1;
	10848 : 1;
	10849 : 1;
	10850 : 1;
	10851 : 1;
	10852 : 1;
	10853 : 1;
	10854 : 1;
	10855 : 1;
	10856 : 1;
	10857 : 1;
	10858 : 1;
	10859 : 1;
	10860 : 1;
	10861 : 1;
	10862 : 1;
	10863 : 1;
	10864 : 1;
	10865 : 1;
	10866 : 1;
	10867 : 1;
	10868 : 1;
	10869 : 1;
	10870 : 1;
	10871 : 1;
	10872 : 1;
	10873 : 1;
	10874 : 1;
	10875 : 1;
	10876 : 1;
	10877 : 1;
	10878 : 1;
	10879 : 1;
	10880 : 1;
	10881 : 1;
	10882 : 1;
	10883 : 1;
	10884 : 1;
	10885 : 1;
	10886 : 1;
	10887 : 1;
	10888 : 1;
	10889 : 1;
	10890 : 1;
	10891 : 1;
	10892 : 1;
	10893 : 1;
	10894 : 1;
	10895 : 1;
	10896 : 1;
	10897 : 1;
	10898 : 1;
	10899 : 1;
	10900 : 1;
	10901 : 1;
	10902 : 1;
	10903 : 1;
	10904 : 1;
	10905 : 1;
	10906 : 1;
	10907 : 1;
	10908 : 1;
	10909 : 1;
	10910 : 1;
	10911 : 1;
	10912 : 1;
	10913 : 1;
	10914 : 1;
	10915 : 1;
	10916 : 1;
	10917 : 1;
	10918 : 1;
	10919 : 1;
	10920 : 1;
	10921 : 1;
	10922 : 1;
	10923 : 1;
	10924 : 1;
	10925 : 1;
	10926 : 1;
	10927 : 1;
	10928 : 1;
	10929 : 1;
	10930 : 1;
	10931 : 1;
	10932 : 1;
	10933 : 1;
	10934 : 1;
	10935 : 1;
	10936 : 1;
	10937 : 1;
	10938 : 1;
	10939 : 1;
	10940 : 1;
	10941 : 1;
	10942 : 1;
	10943 : 1;
	10944 : 1;
	10945 : 1;
	10946 : 1;
	10947 : 1;
	10948 : 1;
	10949 : 1;
	10950 : 1;
	10951 : 1;
	10952 : 1;
	10953 : 1;
	10954 : 1;
	10955 : 1;
	10956 : 1;
	10957 : 1;
	10958 : 1;
	10959 : 1;
	10960 : 1;
	10961 : 1;
	10962 : 1;
	10963 : 1;
	10964 : 1;
	10965 : 1;
	10966 : 1;
	10967 : 1;
	10968 : 1;
	10969 : 1;
	10970 : 1;
	10971 : 1;
	10972 : 1;
	10973 : 1;
	10974 : 1;
	10975 : 1;
	10976 : 1;
	10977 : 1;
	10978 : 1;
	10979 : 1;
	10980 : 1;
	10981 : 1;
	10982 : 1;
	10983 : 1;
	10984 : 1;
	10985 : 1;
	10986 : 1;
	10987 : 1;
	10988 : 1;
	10989 : 1;
	10990 : 1;
	10991 : 1;
	10992 : 1;
	10993 : 1;
	10994 : 1;
	10995 : 1;
	10996 : 1;
	10997 : 1;
	10998 : 1;
	10999 : 1;
	11000 : 1;
	11001 : 1;
	11002 : 1;
	11003 : 1;
	11004 : 1;
	11005 : 1;
	11006 : 1;
	11007 : 1;
	11008 : 1;
	11009 : 1;
	11010 : 1;
	11011 : 1;
	11012 : 1;
	11013 : 1;
	11014 : 1;
	11015 : 1;
	11016 : 1;
	11017 : 1;
	11018 : 1;
	11019 : 1;
	11020 : 1;
	11021 : 1;
	11022 : 1;
	11023 : 1;
	11024 : 1;
	11025 : 1;
	11026 : 1;
	11027 : 1;
	11028 : 1;
	11029 : 1;
	11030 : 1;
	11031 : 1;
	11032 : 1;
	11033 : 1;
	11034 : 1;
	11035 : 1;
	11036 : 1;
	11037 : 1;
	11038 : 1;
	11039 : 1;
	11040 : 1;
	11041 : 1;
	11042 : 1;
	11043 : 1;
	11044 : 1;
	11045 : 1;
	11046 : 1;
	11047 : 1;
	11048 : 1;
	11049 : 1;
	11050 : 1;
	11051 : 1;
	11052 : 1;
	11053 : 1;
	11054 : 1;
	11055 : 1;
	11056 : 1;
	11057 : 1;
	11058 : 1;
	11059 : 1;
	11060 : 1;
	11061 : 1;
	11062 : 1;
	11063 : 1;
	11064 : 1;
	11065 : 1;
	11066 : 1;
	11067 : 1;
	11068 : 1;
	11069 : 1;
	11070 : 1;
	11071 : 1;
	11072 : 1;
	11073 : 1;
	11074 : 1;
	11075 : 1;
	11076 : 1;
	11077 : 1;
	11078 : 1;
	11079 : 1;
	11080 : 1;
	11081 : 1;
	11082 : 1;
	11083 : 1;
	11084 : 1;
	11085 : 1;
	11086 : 1;
	11087 : 1;
	11088 : 1;
	11089 : 1;
	11090 : 1;
	11091 : 1;
	11092 : 1;
	11093 : 1;
	11094 : 1;
	11095 : 1;
	11096 : 1;
	11097 : 1;
	11098 : 1;
	11099 : 1;
	11100 : 1;
	11101 : 1;
	11102 : 1;
	11103 : 1;
	11104 : 1;
	11105 : 1;
	11106 : 1;
	11107 : 1;
	11108 : 1;
	11109 : 1;
	11110 : 1;
	11111 : 1;
	11112 : 1;
	11113 : 1;
	11114 : 1;
	11115 : 1;
	11116 : 1;
	11117 : 1;
	11118 : 1;
	11119 : 1;
	11120 : 1;
	11121 : 1;
	11122 : 1;
	11123 : 1;
	11124 : 1;
	11125 : 1;
	11126 : 1;
	11127 : 1;
	11128 : 1;
	11129 : 1;
	11130 : 1;
	11131 : 1;
	11132 : 1;
	11133 : 1;
	11134 : 1;
	11135 : 1;
	11136 : 1;
	11137 : 1;
	11138 : 1;
	11139 : 1;
	11140 : 1;
	11141 : 1;
	11142 : 1;
	11143 : 1;
	11144 : 1;
	11145 : 1;
	11146 : 1;
	11147 : 1;
	11148 : 1;
	11149 : 1;
	11150 : 1;
	11151 : 1;
	11152 : 1;
	11153 : 1;
	11154 : 1;
	11155 : 1;
	11156 : 1;
	11157 : 1;
	11158 : 1;
	11159 : 1;
	11160 : 1;
	11161 : 1;
	11162 : 1;
	11163 : 1;
	11164 : 1;
	11165 : 1;
	11166 : 1;
	11167 : 1;
	11168 : 1;
	11169 : 1;
	11170 : 1;
	11171 : 1;
	11172 : 1;
	11173 : 1;
	11174 : 1;
	11175 : 1;
	11176 : 1;
	11177 : 1;
	11178 : 1;
	11179 : 1;
	11180 : 1;
	11181 : 1;
	11182 : 1;
	11183 : 1;
	11184 : 1;
	11185 : 1;
	11186 : 1;
	11187 : 1;
	11188 : 1;
	11189 : 1;
	11190 : 1;
	11191 : 1;
	11192 : 1;
	11193 : 1;
	11194 : 1;
	11195 : 1;
	11196 : 1;
	11197 : 1;
	11198 : 1;
	11199 : 1;
	11200 : 1;
	11201 : 1;
	11202 : 1;
	11203 : 1;
	11204 : 1;
	11205 : 1;
	11206 : 1;
	11207 : 1;
	11208 : 1;
	11209 : 1;
	11210 : 1;
	11211 : 1;
	11212 : 1;
	11213 : 1;
	11214 : 1;
	11215 : 1;
	11216 : 1;
	11217 : 1;
	11218 : 1;
	11219 : 1;
	11220 : 1;
	11221 : 1;
	11222 : 1;
	11223 : 1;
	11224 : 1;
	11225 : 1;
	11226 : 1;
	11227 : 1;
	11228 : 1;
	11229 : 1;
	11230 : 1;
	11231 : 1;
	11232 : 1;
	11233 : 1;
	11234 : 1;
	11235 : 1;
	11236 : 1;
	11237 : 1;
	11238 : 1;
	11239 : 1;
	11240 : 1;
	11241 : 1;
	11242 : 1;
	11243 : 1;
	11244 : 1;
	11245 : 1;
	11246 : 1;
	11247 : 1;
	11248 : 1;
	11249 : 1;
	11250 : 1;
	11251 : 1;
	11252 : 1;
	11253 : 1;
	11254 : 1;
	11255 : 1;
	11256 : 1;
	11257 : 1;
	11258 : 1;
	11259 : 1;
	11260 : 1;
	11261 : 1;
	11262 : 1;
	11263 : 1;
	11264 : 1;
	11265 : 1;
	11266 : 1;
	11267 : 1;
	11268 : 1;
	11269 : 1;
	11270 : 1;
	11271 : 1;
	11272 : 1;
	11273 : 1;
	11274 : 1;
	11275 : 1;
	11276 : 1;
	11277 : 1;
	11278 : 1;
	11279 : 1;
	11280 : 1;
	11281 : 1;
	11282 : 1;
	11283 : 1;
	11284 : 1;
	11285 : 1;
	11286 : 1;
	11287 : 1;
	11288 : 1;
	11289 : 1;
	11290 : 1;
	11291 : 1;
	11292 : 1;
	11293 : 1;
	11294 : 1;
	11295 : 1;
	11296 : 1;
	11297 : 1;
	11298 : 1;
	11299 : 1;
	11300 : 1;
	11301 : 1;
	11302 : 1;
	11303 : 1;
	11304 : 1;
	11305 : 1;
	11306 : 1;
	11307 : 1;
	11308 : 1;
	11309 : 1;
	11310 : 1;
	11311 : 1;
	11312 : 1;
	11313 : 1;
	11314 : 1;
	11315 : 1;
	11316 : 1;
	11317 : 1;
	11318 : 1;
	11319 : 1;
	11320 : 1;
	11321 : 1;
	11322 : 1;
	11323 : 1;
	11324 : 1;
	11325 : 1;
	11326 : 1;
	11327 : 1;
	11328 : 1;
	11329 : 1;
	11330 : 1;
	11331 : 1;
	11332 : 1;
	11333 : 1;
	11334 : 1;
	11335 : 1;
	11336 : 1;
	11337 : 1;
	11338 : 1;
	11339 : 1;
	11340 : 1;
	11341 : 1;
	11342 : 1;
	11343 : 1;
	11344 : 1;
	11345 : 1;
	11346 : 1;
	11347 : 1;
	11348 : 1;
	11349 : 1;
	11350 : 1;
	11351 : 1;
	11352 : 1;
	11353 : 1;
	11354 : 1;
	11355 : 1;
	11356 : 1;
	11357 : 1;
	11358 : 1;
	11359 : 1;
	11360 : 1;
	11361 : 1;
	11362 : 1;
	11363 : 1;
	11364 : 1;
	11365 : 1;
	11366 : 1;
	11367 : 1;
	11368 : 1;
	11369 : 1;
	11370 : 1;
	11371 : 1;
	11372 : 1;
	11373 : 1;
	11374 : 1;
	11375 : 1;
	11376 : 1;
	11377 : 1;
	11378 : 1;
	11379 : 1;
	11380 : 1;
	11381 : 1;
	11382 : 1;
	11383 : 1;
	11384 : 1;
	11385 : 1;
	11386 : 1;
	11387 : 1;
	11388 : 1;
	11389 : 1;
	11390 : 1;
	11391 : 1;
	11392 : 1;
	11393 : 1;
	11394 : 1;
	11395 : 1;
	11396 : 1;
	11397 : 1;
	11398 : 1;
	11399 : 1;
	11400 : 1;
	11401 : 1;
	11402 : 1;
	11403 : 1;
	11404 : 1;
	11405 : 1;
	11406 : 1;
	11407 : 1;
	11408 : 1;
	11409 : 1;
	11410 : 1;
	11411 : 1;
	11412 : 1;
	11413 : 1;
	11414 : 1;
	11415 : 1;
	11416 : 1;
	11417 : 1;
	11418 : 1;
	11419 : 1;
	11420 : 1;
	11421 : 1;
	11422 : 1;
	11423 : 1;
	11424 : 1;
	11425 : 1;
	11426 : 1;
	11427 : 1;
	11428 : 1;
	11429 : 1;
	11430 : 1;
	11431 : 1;
	11432 : 1;
	11433 : 1;
	11434 : 1;
	11435 : 1;
	11436 : 1;
	11437 : 1;
	11438 : 1;
	11439 : 1;
	11440 : 1;
	11441 : 1;
	11442 : 1;
	11443 : 1;
	11444 : 1;
	11445 : 1;
	11446 : 1;
	11447 : 1;
	11448 : 1;
	11449 : 1;
	11450 : 1;
	11451 : 1;
	11452 : 1;
	11453 : 1;
	11454 : 1;
	11455 : 1;
	11456 : 1;
	11457 : 1;
	11458 : 1;
	11459 : 1;
	11460 : 1;
	11461 : 1;
	11462 : 1;
	11463 : 1;
	11464 : 1;
	11465 : 1;
	11466 : 1;
	11467 : 1;
	11468 : 1;
	11469 : 1;
	11470 : 1;
	11471 : 1;
	11472 : 1;
	11473 : 1;
	11474 : 1;
	11475 : 1;
	11476 : 1;
	11477 : 1;
	11478 : 1;
	11479 : 1;
	11480 : 1;
	11481 : 1;
	11482 : 1;
	11483 : 1;
	11484 : 1;
	11485 : 1;
	11486 : 1;
	11487 : 1;
	11488 : 1;
	11489 : 1;
	11490 : 1;
	11491 : 1;
	11492 : 1;
	11493 : 1;
	11494 : 1;
	11495 : 1;
	11496 : 1;
	11497 : 1;
	11498 : 1;
	11499 : 1;
	11500 : 1;
	11501 : 1;
	11502 : 1;
	11503 : 1;
	11504 : 1;
	11505 : 1;
	11506 : 1;
	11507 : 1;
	11508 : 1;
	11509 : 1;
	11510 : 1;
	11511 : 1;
	11512 : 1;
	11513 : 1;
	11514 : 1;
	11515 : 1;
	11516 : 1;
	11517 : 1;
	11518 : 1;
	11519 : 1;
	11520 : 1;
	11521 : 1;
	11522 : 1;
	11523 : 1;
	11524 : 1;
	11525 : 1;
	11526 : 1;
	11527 : 1;
	11528 : 1;
	11529 : 1;
	11530 : 1;
	11531 : 1;
	11532 : 1;
	11533 : 1;
	11534 : 1;
	11535 : 1;
	11536 : 1;
	11537 : 1;
	11538 : 1;
	11539 : 1;
	11540 : 1;
	11541 : 1;
	11542 : 1;
	11543 : 1;
	11544 : 1;
	11545 : 1;
	11546 : 1;
	11547 : 1;
	11548 : 1;
	11549 : 1;
	11550 : 1;
	11551 : 1;
	11552 : 1;
	11553 : 1;
	11554 : 1;
	11555 : 1;
	11556 : 1;
	11557 : 1;
	11558 : 1;
	11559 : 1;
	11560 : 1;
	11561 : 1;
	11562 : 1;
	11563 : 1;
	11564 : 1;
	11565 : 1;
	11566 : 1;
	11567 : 1;
	11568 : 1;
	11569 : 1;
	11570 : 1;
	11571 : 1;
	11572 : 1;
	11573 : 1;
	11574 : 1;
	11575 : 1;
	11576 : 1;
	11577 : 1;
	11578 : 1;
	11579 : 1;
	11580 : 1;
	11581 : 1;
	11582 : 1;
	11583 : 1;
	11584 : 1;
	11585 : 1;
	11586 : 1;
	11587 : 1;
	11588 : 1;
	11589 : 1;
	11590 : 1;
	11591 : 1;
	11592 : 1;
	11593 : 1;
	11594 : 1;
	11595 : 1;
	11596 : 1;
	11597 : 1;
	11598 : 1;
	11599 : 1;
	11600 : 1;
	11601 : 1;
	11602 : 1;
	11603 : 1;
	11604 : 1;
	11605 : 1;
	11606 : 1;
	11607 : 1;
	11608 : 1;
	11609 : 1;
	11610 : 1;
	11611 : 1;
	11612 : 1;
	11613 : 1;
	11614 : 1;
	11615 : 1;
	11616 : 1;
	11617 : 1;
	11618 : 1;
	11619 : 1;
	11620 : 1;
	11621 : 1;
	11622 : 1;
	11623 : 1;
	11624 : 1;
	11625 : 1;
	11626 : 1;
	11627 : 1;
	11628 : 1;
	11629 : 1;
	11630 : 1;
	11631 : 1;
	11632 : 1;
	11633 : 1;
	11634 : 1;
	11635 : 1;
	11636 : 1;
	11637 : 1;
	11638 : 1;
	11639 : 1;
	11640 : 1;
	11641 : 1;
	11642 : 1;
	11643 : 1;
	11644 : 1;
	11645 : 1;
	11646 : 1;
	11647 : 1;
	11648 : 1;
	11649 : 1;
	11650 : 1;
	11651 : 1;
	11652 : 1;
	11653 : 1;
	11654 : 1;
	11655 : 1;
	11656 : 1;
	11657 : 1;
	11658 : 1;
	11659 : 1;
	11660 : 1;
	11661 : 1;
	11662 : 1;
	11663 : 1;
	11664 : 1;
	11665 : 1;
	11666 : 1;
	11667 : 1;
	11668 : 1;
	11669 : 1;
	11670 : 1;
	11671 : 1;
	11672 : 1;
	11673 : 1;
	11674 : 1;
	11675 : 1;
	11676 : 1;
	11677 : 1;
	11678 : 1;
	11679 : 1;
	11680 : 1;
	11681 : 1;
	11682 : 1;
	11683 : 1;
	11684 : 1;
	11685 : 1;
	11686 : 1;
	11687 : 1;
	11688 : 1;
	11689 : 1;
	11690 : 1;
	11691 : 1;
	11692 : 1;
	11693 : 1;
	11694 : 1;
	11695 : 1;
	11696 : 1;
	11697 : 1;
	11698 : 1;
	11699 : 1;
	11700 : 1;
	11701 : 1;
	11702 : 1;
	11703 : 1;
	11704 : 1;
	11705 : 1;
	11706 : 1;
	11707 : 1;
	11708 : 1;
	11709 : 1;
	11710 : 1;
	11711 : 1;
	11712 : 1;
	11713 : 1;
	11714 : 1;
	11715 : 1;
	11716 : 1;
	11717 : 1;
	11718 : 1;
	11719 : 1;
	11720 : 1;
	11721 : 1;
	11722 : 1;
	11723 : 1;
	11724 : 1;
	11725 : 1;
	11726 : 1;
	11727 : 1;
	11728 : 1;
	11729 : 1;
	11730 : 1;
	11731 : 1;
	11732 : 1;
	11733 : 1;
	11734 : 1;
	11735 : 1;
	11736 : 1;
	11737 : 1;
	11738 : 1;
	11739 : 1;
	11740 : 1;
	11741 : 1;
	11742 : 1;
	11743 : 1;
	11744 : 1;
	11745 : 1;
	11746 : 1;
	11747 : 1;
	11748 : 1;
	11749 : 1;
	11750 : 1;
	11751 : 1;
	11752 : 1;
	11753 : 1;
	11754 : 1;
	11755 : 1;
	11756 : 1;
	11757 : 1;
	11758 : 1;
	11759 : 1;
	11760 : 1;
	11761 : 1;
	11762 : 1;
	11763 : 1;
	11764 : 1;
	11765 : 1;
	11766 : 1;
	11767 : 1;
	11768 : 1;
	11769 : 1;
	11770 : 1;
	11771 : 1;
	11772 : 1;
	11773 : 1;
	11774 : 1;
	11775 : 1;
	11776 : 1;
	11777 : 1;
	11778 : 1;
	11779 : 1;
	11780 : 1;
	11781 : 1;
	11782 : 1;
	11783 : 1;
	11784 : 1;
	11785 : 1;
	11786 : 1;
	11787 : 1;
	11788 : 1;
	11789 : 1;
	11790 : 1;
	11791 : 1;
	11792 : 1;
	11793 : 1;
	11794 : 1;
	11795 : 1;
	11796 : 1;
	11797 : 1;
	11798 : 1;
	11799 : 1;
	11800 : 1;
	11801 : 1;
	11802 : 1;
	11803 : 1;
	11804 : 1;
	11805 : 1;
	11806 : 1;
	11807 : 1;
	11808 : 1;
	11809 : 1;
	11810 : 1;
	11811 : 1;
	11812 : 1;
	11813 : 1;
	11814 : 1;
	11815 : 1;
	11816 : 1;
	11817 : 1;
	11818 : 1;
	11819 : 1;
	11820 : 1;
	11821 : 1;
	11822 : 1;
	11823 : 1;
	11824 : 1;
	11825 : 1;
	11826 : 1;
	11827 : 1;
	11828 : 1;
	11829 : 1;
	11830 : 1;
	11831 : 1;
	11832 : 1;
	11833 : 1;
	11834 : 1;
	11835 : 1;
	11836 : 1;
	11837 : 1;
	11838 : 1;
	11839 : 1;
	11840 : 1;
	11841 : 1;
	11842 : 1;
	11843 : 1;
	11844 : 1;
	11845 : 1;
	11846 : 1;
	11847 : 1;
	11848 : 1;
	11849 : 1;
	11850 : 1;
	11851 : 1;
	11852 : 1;
	11853 : 1;
	11854 : 1;
	11855 : 1;
	11856 : 1;
	11857 : 1;
	11858 : 1;
	11859 : 1;
	11860 : 1;
	11861 : 1;
	11862 : 1;
	11863 : 1;
	11864 : 1;
	11865 : 1;
	11866 : 1;
	11867 : 1;
	11868 : 1;
	11869 : 1;
	11870 : 1;
	11871 : 1;
	11872 : 1;
	11873 : 1;
	11874 : 1;
	11875 : 1;
	11876 : 1;
	11877 : 1;
	11878 : 1;
	11879 : 1;
	11880 : 1;
	11881 : 1;
	11882 : 1;
	11883 : 1;
	11884 : 1;
	11885 : 1;
	11886 : 1;
	11887 : 1;
	11888 : 1;
	11889 : 1;
	11890 : 1;
	11891 : 1;
	11892 : 1;
	11893 : 1;
	11894 : 1;
	11895 : 1;
	11896 : 1;
	11897 : 1;
	11898 : 1;
	11899 : 1;
	11900 : 1;
	11901 : 1;
	11902 : 1;
	11903 : 1;
	11904 : 1;
	11905 : 1;
	11906 : 1;
	11907 : 1;
	11908 : 1;
	11909 : 1;
	11910 : 1;
	11911 : 1;
	11912 : 1;
	11913 : 1;
	11914 : 1;
	11915 : 1;
	11916 : 1;
	11917 : 1;
	11918 : 1;
	11919 : 1;
	11920 : 1;
	11921 : 1;
	11922 : 1;
	11923 : 1;
	11924 : 1;
	11925 : 1;
	11926 : 1;
	11927 : 1;
	11928 : 1;
	11929 : 1;
	11930 : 1;
	11931 : 1;
	11932 : 1;
	11933 : 1;
	11934 : 1;
	11935 : 1;
	11936 : 1;
	11937 : 1;
	11938 : 1;
	11939 : 1;
	11940 : 1;
	11941 : 1;
	11942 : 1;
	11943 : 1;
	11944 : 1;
	11945 : 1;
	11946 : 1;
	11947 : 1;
	11948 : 1;
	11949 : 1;
	11950 : 1;
	11951 : 1;
	11952 : 1;
	11953 : 1;
	11954 : 1;
	11955 : 1;
	11956 : 1;
	11957 : 1;
	11958 : 1;
	11959 : 1;
	11960 : 1;
	11961 : 1;
	11962 : 1;
	11963 : 1;
	11964 : 1;
	11965 : 1;
	11966 : 1;
	11967 : 1;
	11968 : 1;
	11969 : 1;
	11970 : 1;
	11971 : 1;
	11972 : 1;
	11973 : 1;
	11974 : 1;
	11975 : 1;
	11976 : 1;
	11977 : 1;
	11978 : 1;
	11979 : 1;
	11980 : 1;
	11981 : 1;
	11982 : 1;
	11983 : 1;
	11984 : 1;
	11985 : 1;
	11986 : 1;
	11987 : 1;
	11988 : 1;
	11989 : 1;
	11990 : 1;
	11991 : 1;
	11992 : 1;
	11993 : 1;
	11994 : 1;
	11995 : 1;
	11996 : 1;
	11997 : 1;
	11998 : 1;
	11999 : 1;
	12000 : 1;
	12001 : 1;
	12002 : 1;
	12003 : 1;
	12004 : 1;
	12005 : 1;
	12006 : 1;
	12007 : 1;
	12008 : 1;
	12009 : 1;
	12010 : 1;
	12011 : 1;
	12012 : 1;
	12013 : 1;
	12014 : 1;
	12015 : 1;
	12016 : 1;
	12017 : 1;
	12018 : 1;
	12019 : 1;
	12020 : 1;
	12021 : 1;
	12022 : 1;
	12023 : 1;
	12024 : 1;
	12025 : 1;
	12026 : 1;
	12027 : 1;
	12028 : 1;
	12029 : 1;
	12030 : 1;
	12031 : 1;
	12032 : 1;
	12033 : 1;
	12034 : 1;
	12035 : 1;
	12036 : 1;
	12037 : 1;
	12038 : 1;
	12039 : 1;
	12040 : 1;
	12041 : 1;
	12042 : 1;
	12043 : 1;
	12044 : 1;
	12045 : 1;
	12046 : 1;
	12047 : 1;
	12048 : 1;
	12049 : 1;
	12050 : 1;
	12051 : 1;
	12052 : 1;
	12053 : 1;
	12054 : 1;
	12055 : 1;
	12056 : 1;
	12057 : 1;
	12058 : 1;
	12059 : 1;
	12060 : 1;
	12061 : 1;
	12062 : 1;
	12063 : 1;
	12064 : 1;
	12065 : 1;
	12066 : 1;
	12067 : 1;
	12068 : 1;
	12069 : 1;
	12070 : 1;
	12071 : 1;
	12072 : 1;
	12073 : 1;
	12074 : 1;
	12075 : 1;
	12076 : 1;
	12077 : 1;
	12078 : 1;
	12079 : 1;
	12080 : 1;
	12081 : 1;
	12082 : 1;
	12083 : 1;
	12084 : 1;
	12085 : 1;
	12086 : 1;
	12087 : 1;
	12088 : 1;
	12089 : 1;
	12090 : 1;
	12091 : 1;
	12092 : 1;
	12093 : 1;
	12094 : 1;
	12095 : 1;
	12096 : 1;
	12097 : 1;
	12098 : 1;
	12099 : 1;
	12100 : 1;
	12101 : 1;
	12102 : 1;
	12103 : 1;
	12104 : 1;
	12105 : 1;
	12106 : 1;
	12107 : 1;
	12108 : 1;
	12109 : 1;
	12110 : 1;
	12111 : 1;
	12112 : 1;
	12113 : 1;
	12114 : 1;
	12115 : 1;
	12116 : 1;
	12117 : 1;
	12118 : 1;
	12119 : 1;
	12120 : 1;
	12121 : 1;
	12122 : 1;
	12123 : 1;
	12124 : 1;
	12125 : 1;
	12126 : 1;
	12127 : 1;
	12128 : 1;
	12129 : 1;
	12130 : 1;
	12131 : 1;
	12132 : 1;
	12133 : 1;
	12134 : 1;
	12135 : 1;
	12136 : 1;
	12137 : 1;
	12138 : 1;
	12139 : 1;
	12140 : 1;
	12141 : 1;
	12142 : 1;
	12143 : 1;
	12144 : 1;
	12145 : 1;
	12146 : 1;
	12147 : 1;
	12148 : 1;
	12149 : 1;
	12150 : 1;
	12151 : 1;
	12152 : 1;
	12153 : 1;
	12154 : 1;
	12155 : 1;
	12156 : 1;
	12157 : 1;
	12158 : 1;
	12159 : 1;
	12160 : 1;
	12161 : 1;
	12162 : 1;
	12163 : 1;
	12164 : 1;
	12165 : 1;
	12166 : 1;
	12167 : 1;
	12168 : 1;
	12169 : 1;
	12170 : 1;
	12171 : 1;
	12172 : 1;
	12173 : 1;
	12174 : 1;
	12175 : 1;
	12176 : 1;
	12177 : 1;
	12178 : 1;
	12179 : 1;
	12180 : 1;
	12181 : 1;
	12182 : 1;
	12183 : 1;
	12184 : 1;
	12185 : 1;
	12186 : 1;
	12187 : 1;
	12188 : 1;
	12189 : 1;
	12190 : 1;
	12191 : 1;
	12192 : 1;
	12193 : 1;
	12194 : 1;
	12195 : 1;
	12196 : 1;
	12197 : 1;
	12198 : 1;
	12199 : 1;
	12200 : 1;
	12201 : 1;
	12202 : 1;
	12203 : 1;
	12204 : 1;
	12205 : 1;
	12206 : 1;
	12207 : 1;
	12208 : 1;
	12209 : 1;
	12210 : 1;
	12211 : 1;
	12212 : 1;
	12213 : 1;
	12214 : 1;
	12215 : 1;
	12216 : 1;
	12217 : 1;
	12218 : 1;
	12219 : 1;
	12220 : 1;
	12221 : 1;
	12222 : 1;
	12223 : 1;
	12224 : 1;
	12225 : 1;
	12226 : 1;
	12227 : 1;
	12228 : 1;
	12229 : 1;
	12230 : 1;
	12231 : 1;
	12232 : 1;
	12233 : 1;
	12234 : 1;
	12235 : 1;
	12236 : 1;
	12237 : 1;
	12238 : 1;
	12239 : 1;
	12240 : 1;
	12241 : 1;
	12242 : 1;
	12243 : 1;
	12244 : 1;
	12245 : 1;
	12246 : 1;
	12247 : 1;
	12248 : 1;
	12249 : 1;
	12250 : 1;
	12251 : 1;
	12252 : 1;
	12253 : 1;
	12254 : 1;
	12255 : 1;
	12256 : 1;
	12257 : 1;
	12258 : 1;
	12259 : 1;
	12260 : 1;
	12261 : 1;
	12262 : 1;
	12263 : 1;
	12264 : 1;
	12265 : 1;
	12266 : 1;
	12267 : 1;
	12268 : 1;
	12269 : 1;
	12270 : 0;
	12271 : 0;
	12272 : 0;
	12273 : 0;
	12274 : 1;
	12275 : 1;
	12276 : 1;
	12277 : 1;
	12278 : 1;
	12279 : 1;
	12280 : 1;
	12281 : 1;
	12282 : 1;
	12283 : 1;
	12284 : 1;
	12285 : 1;
	12286 : 1;
	12287 : 1;
	12288 : 1;
	12289 : 1;
	12290 : 1;
	12291 : 1;
	12292 : 1;
	12293 : 1;
	12294 : 0;
	12295 : 1;
	12296 : 1;
	12297 : 1;
	12298 : 1;
	12299 : 1;
	12300 : 1;
	12301 : 1;
	12302 : 1;
	12303 : 0;
	12304 : 0;
	12305 : 1;
	12306 : 1;
	12307 : 1;
	12308 : 1;
	12309 : 1;
	12310 : 1;
	12311 : 1;
	12312 : 1;
	12313 : 0;
	12314 : 1;
	12315 : 1;
	12316 : 1;
	12317 : 1;
	12318 : 1;
	12319 : 1;
	12320 : 1;
	12321 : 1;
	12322 : 1;
	12323 : 1;
	12324 : 1;
	12325 : 1;
	12326 : 1;
	12327 : 1;
	12328 : 1;
	12329 : 1;
	12330 : 1;
	12331 : 0;
	12332 : 1;
	12333 : 1;
	12334 : 1;
	12335 : 1;
	12336 : 1;
	12337 : 1;
	12338 : 1;
	12339 : 1;
	12340 : 1;
	12341 : 1;
	12342 : 1;
	12343 : 1;
	12344 : 1;
	12345 : 1;
	12346 : 1;
	12347 : 1;
	12348 : 1;
	12349 : 1;
	12350 : 1;
	12351 : 1;
	12352 : 1;
	12353 : 1;
	12354 : 1;
	12355 : 1;
	12356 : 1;
	12357 : 1;
	12358 : 1;
	12359 : 1;
	12360 : 1;
	12361 : 1;
	12362 : 1;
	12363 : 1;
	12364 : 1;
	12365 : 1;
	12366 : 1;
	12367 : 1;
	12368 : 1;
	12369 : 1;
	12370 : 1;
	12371 : 1;
	12372 : 1;
	12373 : 1;
	12374 : 1;
	12375 : 1;
	12376 : 1;
	12377 : 0;
	12378 : 0;
	12379 : 0;
	12380 : 0;
	12381 : 0;
	12382 : 1;
	12383 : 0;
	12384 : 0;
	12385 : 0;
	12386 : 0;
	12387 : 1;
	12388 : 1;
	12389 : 1;
	12390 : 1;
	12391 : 0;
	12392 : 0;
	12393 : 0;
	12394 : 0;
	12395 : 0;
	12396 : 1;
	12397 : 1;
	12398 : 1;
	12399 : 1;
	12400 : 1;
	12401 : 1;
	12402 : 1;
	12403 : 0;
	12404 : 0;
	12405 : 1;
	12406 : 1;
	12407 : 1;
	12408 : 1;
	12409 : 1;
	12410 : 1;
	12411 : 1;
	12412 : 1;
	12413 : 1;
	12414 : 1;
	12415 : 1;
	12416 : 1;
	12417 : 1;
	12418 : 1;
	12419 : 1;
	12420 : 1;
	12421 : 1;
	12422 : 1;
	12423 : 1;
	12424 : 1;
	12425 : 1;
	12426 : 1;
	12427 : 0;
	12428 : 0;
	12429 : 1;
	12430 : 1;
	12431 : 1;
	12432 : 1;
	12433 : 1;
	12434 : 1;
	12435 : 1;
	12436 : 1;
	12437 : 1;
	12438 : 1;
	12439 : 1;
	12440 : 1;
	12441 : 1;
	12442 : 1;
	12443 : 1;
	12444 : 1;
	12445 : 1;
	12446 : 1;
	12447 : 1;
	12448 : 1;
	12449 : 1;
	12450 : 1;
	12451 : 1;
	12452 : 1;
	12453 : 1;
	12454 : 1;
	12455 : 1;
	12456 : 1;
	12457 : 1;
	12458 : 1;
	12459 : 1;
	12460 : 1;
	12461 : 1;
	12462 : 1;
	12463 : 1;
	12464 : 1;
	12465 : 1;
	12466 : 1;
	12467 : 1;
	12468 : 1;
	12469 : 1;
	12470 : 1;
	12471 : 1;
	12472 : 1;
	12473 : 1;
	12474 : 1;
	12475 : 1;
	12476 : 1;
	12477 : 1;
	12478 : 1;
	12479 : 1;
	12480 : 1;
	12481 : 1;
	12482 : 1;
	12483 : 1;
	12484 : 1;
	12485 : 1;
	12486 : 1;
	12487 : 1;
	12488 : 1;
	12489 : 1;
	12490 : 1;
	12491 : 1;
	12492 : 1;
	12493 : 1;
	12494 : 1;
	12495 : 1;
	12496 : 1;
	12497 : 1;
	12498 : 1;
	12499 : 1;
	12500 : 1;
	12501 : 1;
	12502 : 1;
	12503 : 1;
	12504 : 1;
	12505 : 1;
	12506 : 1;
	12507 : 1;
	12508 : 1;
	12509 : 0;
	12510 : 1;
	12511 : 1;
	12512 : 1;
	12513 : 1;
	12514 : 1;
	12515 : 1;
	12516 : 1;
	12517 : 1;
	12518 : 1;
	12519 : 1;
	12520 : 1;
	12521 : 1;
	12522 : 1;
	12523 : 1;
	12524 : 1;
	12525 : 1;
	12526 : 1;
	12527 : 1;
	12528 : 1;
	12529 : 1;
	12530 : 1;
	12531 : 1;
	12532 : 1;
	12533 : 1;
	12534 : 1;
	12535 : 1;
	12536 : 1;
	12537 : 1;
	12538 : 1;
	12539 : 1;
	12540 : 1;
	12541 : 1;
	12542 : 1;
	12543 : 0;
	12544 : 0;
	12545 : 1;
	12546 : 1;
	12547 : 1;
	12548 : 1;
	12549 : 0;
	12550 : 1;
	12551 : 1;
	12552 : 1;
	12553 : 0;
	12554 : 1;
	12555 : 1;
	12556 : 1;
	12557 : 1;
	12558 : 1;
	12559 : 1;
	12560 : 1;
	12561 : 1;
	12562 : 1;
	12563 : 1;
	12564 : 1;
	12565 : 1;
	12566 : 1;
	12567 : 1;
	12568 : 1;
	12569 : 1;
	12570 : 1;
	12571 : 0;
	12572 : 1;
	12573 : 1;
	12574 : 1;
	12575 : 1;
	12576 : 1;
	12577 : 1;
	12578 : 1;
	12579 : 1;
	12580 : 1;
	12581 : 1;
	12582 : 1;
	12583 : 1;
	12584 : 0;
	12585 : 1;
	12586 : 1;
	12587 : 1;
	12588 : 1;
	12589 : 1;
	12590 : 1;
	12591 : 1;
	12592 : 1;
	12593 : 1;
	12594 : 1;
	12595 : 1;
	12596 : 1;
	12597 : 1;
	12598 : 1;
	12599 : 1;
	12600 : 1;
	12601 : 1;
	12602 : 1;
	12603 : 1;
	12604 : 1;
	12605 : 1;
	12606 : 1;
	12607 : 1;
	12608 : 1;
	12609 : 1;
	12610 : 1;
	12611 : 1;
	12612 : 1;
	12613 : 1;
	12614 : 1;
	12615 : 1;
	12616 : 1;
	12617 : 1;
	12618 : 0;
	12619 : 0;
	12620 : 1;
	12621 : 1;
	12622 : 1;
	12623 : 0;
	12624 : 1;
	12625 : 1;
	12626 : 1;
	12627 : 0;
	12628 : 1;
	12629 : 1;
	12630 : 1;
	12631 : 0;
	12632 : 1;
	12633 : 1;
	12634 : 1;
	12635 : 0;
	12636 : 1;
	12637 : 1;
	12638 : 1;
	12639 : 1;
	12640 : 1;
	12641 : 1;
	12642 : 1;
	12643 : 0;
	12644 : 0;
	12645 : 1;
	12646 : 1;
	12647 : 1;
	12648 : 1;
	12649 : 1;
	12650 : 1;
	12651 : 1;
	12652 : 1;
	12653 : 1;
	12654 : 1;
	12655 : 1;
	12656 : 1;
	12657 : 1;
	12658 : 1;
	12659 : 1;
	12660 : 1;
	12661 : 1;
	12662 : 1;
	12663 : 1;
	12664 : 1;
	12665 : 1;
	12666 : 1;
	12667 : 0;
	12668 : 0;
	12669 : 1;
	12670 : 1;
	12671 : 1;
	12672 : 1;
	12673 : 1;
	12674 : 1;
	12675 : 1;
	12676 : 1;
	12677 : 1;
	12678 : 1;
	12679 : 1;
	12680 : 1;
	12681 : 1;
	12682 : 1;
	12683 : 1;
	12684 : 1;
	12685 : 1;
	12686 : 1;
	12687 : 1;
	12688 : 1;
	12689 : 1;
	12690 : 1;
	12691 : 1;
	12692 : 1;
	12693 : 1;
	12694 : 1;
	12695 : 1;
	12696 : 1;
	12697 : 1;
	12698 : 1;
	12699 : 1;
	12700 : 1;
	12701 : 1;
	12702 : 1;
	12703 : 1;
	12704 : 1;
	12705 : 1;
	12706 : 1;
	12707 : 1;
	12708 : 1;
	12709 : 1;
	12710 : 1;
	12711 : 1;
	12712 : 1;
	12713 : 1;
	12714 : 1;
	12715 : 1;
	12716 : 1;
	12717 : 1;
	12718 : 1;
	12719 : 1;
	12720 : 1;
	12721 : 1;
	12722 : 1;
	12723 : 1;
	12724 : 1;
	12725 : 1;
	12726 : 1;
	12727 : 1;
	12728 : 1;
	12729 : 1;
	12730 : 1;
	12731 : 1;
	12732 : 1;
	12733 : 1;
	12734 : 1;
	12735 : 1;
	12736 : 1;
	12737 : 1;
	12738 : 1;
	12739 : 1;
	12740 : 1;
	12741 : 1;
	12742 : 1;
	12743 : 1;
	12744 : 1;
	12745 : 1;
	12746 : 1;
	12747 : 1;
	12748 : 1;
	12749 : 0;
	12750 : 0;
	12751 : 1;
	12752 : 1;
	12753 : 1;
	12754 : 1;
	12755 : 1;
	12756 : 1;
	12757 : 1;
	12758 : 1;
	12759 : 1;
	12760 : 1;
	12761 : 1;
	12762 : 1;
	12763 : 1;
	12764 : 1;
	12765 : 1;
	12766 : 1;
	12767 : 1;
	12768 : 1;
	12769 : 1;
	12770 : 1;
	12771 : 1;
	12772 : 1;
	12773 : 1;
	12774 : 1;
	12775 : 1;
	12776 : 1;
	12777 : 1;
	12778 : 1;
	12779 : 1;
	12780 : 1;
	12781 : 1;
	12782 : 1;
	12783 : 0;
	12784 : 0;
	12785 : 1;
	12786 : 1;
	12787 : 1;
	12788 : 0;
	12789 : 0;
	12790 : 1;
	12791 : 1;
	12792 : 1;
	12793 : 0;
	12794 : 1;
	12795 : 1;
	12796 : 1;
	12797 : 1;
	12798 : 1;
	12799 : 1;
	12800 : 1;
	12801 : 1;
	12802 : 1;
	12803 : 1;
	12804 : 1;
	12805 : 1;
	12806 : 1;
	12807 : 1;
	12808 : 1;
	12809 : 1;
	12810 : 1;
	12811 : 0;
	12812 : 1;
	12813 : 1;
	12814 : 1;
	12815 : 1;
	12816 : 1;
	12817 : 1;
	12818 : 1;
	12819 : 1;
	12820 : 1;
	12821 : 1;
	12822 : 1;
	12823 : 1;
	12824 : 0;
	12825 : 0;
	12826 : 1;
	12827 : 1;
	12828 : 1;
	12829 : 1;
	12830 : 1;
	12831 : 1;
	12832 : 1;
	12833 : 1;
	12834 : 1;
	12835 : 1;
	12836 : 1;
	12837 : 1;
	12838 : 1;
	12839 : 1;
	12840 : 1;
	12841 : 1;
	12842 : 1;
	12843 : 1;
	12844 : 1;
	12845 : 1;
	12846 : 1;
	12847 : 1;
	12848 : 1;
	12849 : 1;
	12850 : 1;
	12851 : 1;
	12852 : 1;
	12853 : 1;
	12854 : 1;
	12855 : 1;
	12856 : 1;
	12857 : 1;
	12858 : 0;
	12859 : 0;
	12860 : 1;
	12861 : 1;
	12862 : 1;
	12863 : 0;
	12864 : 1;
	12865 : 1;
	12866 : 1;
	12867 : 0;
	12868 : 1;
	12869 : 1;
	12870 : 1;
	12871 : 0;
	12872 : 1;
	12873 : 1;
	12874 : 1;
	12875 : 0;
	12876 : 1;
	12877 : 1;
	12878 : 1;
	12879 : 1;
	12880 : 1;
	12881 : 1;
	12882 : 1;
	12883 : 0;
	12884 : 0;
	12885 : 1;
	12886 : 1;
	12887 : 1;
	12888 : 1;
	12889 : 1;
	12890 : 1;
	12891 : 1;
	12892 : 1;
	12893 : 1;
	12894 : 1;
	12895 : 1;
	12896 : 1;
	12897 : 1;
	12898 : 1;
	12899 : 1;
	12900 : 1;
	12901 : 1;
	12902 : 1;
	12903 : 1;
	12904 : 1;
	12905 : 1;
	12906 : 1;
	12907 : 0;
	12908 : 0;
	12909 : 1;
	12910 : 1;
	12911 : 1;
	12912 : 1;
	12913 : 1;
	12914 : 1;
	12915 : 1;
	12916 : 1;
	12917 : 1;
	12918 : 1;
	12919 : 1;
	12920 : 1;
	12921 : 1;
	12922 : 1;
	12923 : 1;
	12924 : 1;
	12925 : 1;
	12926 : 1;
	12927 : 1;
	12928 : 1;
	12929 : 1;
	12930 : 1;
	12931 : 1;
	12932 : 1;
	12933 : 1;
	12934 : 1;
	12935 : 1;
	12936 : 1;
	12937 : 1;
	12938 : 1;
	12939 : 1;
	12940 : 1;
	12941 : 1;
	12942 : 1;
	12943 : 1;
	12944 : 1;
	12945 : 1;
	12946 : 1;
	12947 : 1;
	12948 : 1;
	12949 : 1;
	12950 : 1;
	12951 : 1;
	12952 : 1;
	12953 : 1;
	12954 : 1;
	12955 : 1;
	12956 : 1;
	12957 : 1;
	12958 : 1;
	12959 : 1;
	12960 : 1;
	12961 : 1;
	12962 : 1;
	12963 : 1;
	12964 : 1;
	12965 : 1;
	12966 : 1;
	12967 : 1;
	12968 : 1;
	12969 : 1;
	12970 : 1;
	12971 : 1;
	12972 : 1;
	12973 : 1;
	12974 : 1;
	12975 : 1;
	12976 : 1;
	12977 : 1;
	12978 : 1;
	12979 : 1;
	12980 : 1;
	12981 : 1;
	12982 : 1;
	12983 : 1;
	12984 : 1;
	12985 : 1;
	12986 : 1;
	12987 : 1;
	12988 : 1;
	12989 : 1;
	12990 : 0;
	12991 : 0;
	12992 : 0;
	12993 : 1;
	12994 : 1;
	12995 : 0;
	12996 : 0;
	12997 : 0;
	12998 : 0;
	12999 : 0;
	13000 : 1;
	13001 : 1;
	13002 : 0;
	13003 : 0;
	13004 : 0;
	13005 : 0;
	13006 : 1;
	13007 : 1;
	13008 : 1;
	13009 : 0;
	13010 : 0;
	13011 : 0;
	13012 : 0;
	13013 : 1;
	13014 : 0;
	13015 : 1;
	13016 : 1;
	13017 : 0;
	13018 : 0;
	13019 : 0;
	13020 : 0;
	13021 : 0;
	13022 : 1;
	13023 : 0;
	13024 : 0;
	13025 : 1;
	13026 : 1;
	13027 : 1;
	13028 : 0;
	13029 : 0;
	13030 : 0;
	13031 : 0;
	13032 : 1;
	13033 : 0;
	13034 : 0;
	13035 : 0;
	13036 : 0;
	13037 : 0;
	13038 : 1;
	13039 : 1;
	13040 : 0;
	13041 : 0;
	13042 : 0;
	13043 : 0;
	13044 : 0;
	13045 : 0;
	13046 : 0;
	13047 : 0;
	13048 : 0;
	13049 : 1;
	13050 : 1;
	13051 : 0;
	13052 : 1;
	13053 : 0;
	13054 : 0;
	13055 : 1;
	13056 : 0;
	13057 : 0;
	13058 : 0;
	13059 : 0;
	13060 : 1;
	13061 : 1;
	13062 : 1;
	13063 : 0;
	13064 : 0;
	13065 : 0;
	13066 : 0;
	13067 : 1;
	13068 : 1;
	13069 : 0;
	13070 : 0;
	13071 : 0;
	13072 : 0;
	13073 : 1;
	13074 : 1;
	13075 : 1;
	13076 : 1;
	13077 : 0;
	13078 : 0;
	13079 : 0;
	13080 : 0;
	13081 : 1;
	13082 : 1;
	13083 : 0;
	13084 : 1;
	13085 : 1;
	13086 : 0;
	13087 : 1;
	13088 : 1;
	13089 : 0;
	13090 : 0;
	13091 : 0;
	13092 : 0;
	13093 : 1;
	13094 : 1;
	13095 : 1;
	13096 : 1;
	13097 : 1;
	13098 : 0;
	13099 : 0;
	13100 : 1;
	13101 : 1;
	13102 : 1;
	13103 : 0;
	13104 : 1;
	13105 : 1;
	13106 : 1;
	13107 : 0;
	13108 : 1;
	13109 : 1;
	13110 : 1;
	13111 : 0;
	13112 : 1;
	13113 : 1;
	13114 : 1;
	13115 : 0;
	13116 : 1;
	13117 : 1;
	13118 : 0;
	13119 : 0;
	13120 : 0;
	13121 : 0;
	13122 : 1;
	13123 : 0;
	13124 : 0;
	13125 : 0;
	13126 : 0;
	13127 : 0;
	13128 : 1;
	13129 : 1;
	13130 : 0;
	13131 : 1;
	13132 : 1;
	13133 : 0;
	13134 : 1;
	13135 : 1;
	13136 : 0;
	13137 : 0;
	13138 : 0;
	13139 : 0;
	13140 : 1;
	13141 : 1;
	13142 : 1;
	13143 : 1;
	13144 : 1;
	13145 : 1;
	13146 : 1;
	13147 : 0;
	13148 : 0;
	13149 : 1;
	13150 : 0;
	13151 : 0;
	13152 : 0;
	13153 : 0;
	13154 : 1;
	13155 : 1;
	13156 : 0;
	13157 : 0;
	13158 : 0;
	13159 : 0;
	13160 : 1;
	13161 : 1;
	13162 : 0;
	13163 : 0;
	13164 : 0;
	13165 : 0;
	13166 : 1;
	13167 : 1;
	13168 : 1;
	13169 : 1;
	13170 : 1;
	13171 : 1;
	13172 : 1;
	13173 : 1;
	13174 : 1;
	13175 : 1;
	13176 : 1;
	13177 : 1;
	13178 : 1;
	13179 : 1;
	13180 : 1;
	13181 : 1;
	13182 : 1;
	13183 : 1;
	13184 : 1;
	13185 : 1;
	13186 : 1;
	13187 : 1;
	13188 : 1;
	13189 : 1;
	13190 : 1;
	13191 : 1;
	13192 : 1;
	13193 : 1;
	13194 : 1;
	13195 : 1;
	13196 : 1;
	13197 : 1;
	13198 : 1;
	13199 : 1;
	13200 : 1;
	13201 : 1;
	13202 : 1;
	13203 : 1;
	13204 : 1;
	13205 : 1;
	13206 : 1;
	13207 : 1;
	13208 : 1;
	13209 : 1;
	13210 : 1;
	13211 : 1;
	13212 : 1;
	13213 : 1;
	13214 : 1;
	13215 : 1;
	13216 : 1;
	13217 : 1;
	13218 : 1;
	13219 : 1;
	13220 : 1;
	13221 : 1;
	13222 : 1;
	13223 : 1;
	13224 : 1;
	13225 : 1;
	13226 : 1;
	13227 : 1;
	13228 : 1;
	13229 : 1;
	13230 : 1;
	13231 : 1;
	13232 : 0;
	13233 : 0;
	13234 : 1;
	13235 : 0;
	13236 : 0;
	13237 : 1;
	13238 : 1;
	13239 : 1;
	13240 : 0;
	13241 : 1;
	13242 : 0;
	13243 : 1;
	13244 : 1;
	13245 : 1;
	13246 : 0;
	13247 : 1;
	13248 : 0;
	13249 : 1;
	13250 : 1;
	13251 : 1;
	13252 : 0;
	13253 : 1;
	13254 : 0;
	13255 : 1;
	13256 : 0;
	13257 : 1;
	13258 : 1;
	13259 : 1;
	13260 : 0;
	13261 : 0;
	13262 : 1;
	13263 : 0;
	13264 : 0;
	13265 : 1;
	13266 : 1;
	13267 : 1;
	13268 : 1;
	13269 : 0;
	13270 : 1;
	13271 : 1;
	13272 : 1;
	13273 : 0;
	13274 : 1;
	13275 : 1;
	13276 : 1;
	13277 : 0;
	13278 : 1;
	13279 : 0;
	13280 : 1;
	13281 : 1;
	13282 : 1;
	13283 : 0;
	13284 : 0;
	13285 : 0;
	13286 : 0;
	13287 : 1;
	13288 : 0;
	13289 : 0;
	13290 : 1;
	13291 : 0;
	13292 : 0;
	13293 : 0;
	13294 : 1;
	13295 : 1;
	13296 : 0;
	13297 : 1;
	13298 : 1;
	13299 : 1;
	13300 : 1;
	13301 : 1;
	13302 : 1;
	13303 : 1;
	13304 : 0;
	13305 : 1;
	13306 : 1;
	13307 : 1;
	13308 : 0;
	13309 : 1;
	13310 : 1;
	13311 : 1;
	13312 : 0;
	13313 : 0;
	13314 : 1;
	13315 : 1;
	13316 : 1;
	13317 : 0;
	13318 : 1;
	13319 : 1;
	13320 : 1;
	13321 : 0;
	13322 : 1;
	13323 : 0;
	13324 : 1;
	13325 : 1;
	13326 : 0;
	13327 : 1;
	13328 : 1;
	13329 : 0;
	13330 : 0;
	13331 : 1;
	13332 : 1;
	13333 : 1;
	13334 : 1;
	13335 : 1;
	13336 : 1;
	13337 : 1;
	13338 : 0;
	13339 : 0;
	13340 : 1;
	13341 : 1;
	13342 : 1;
	13343 : 0;
	13344 : 0;
	13345 : 0;
	13346 : 0;
	13347 : 0;
	13348 : 1;
	13349 : 1;
	13350 : 1;
	13351 : 0;
	13352 : 1;
	13353 : 1;
	13354 : 1;
	13355 : 0;
	13356 : 1;
	13357 : 0;
	13358 : 1;
	13359 : 1;
	13360 : 1;
	13361 : 0;
	13362 : 0;
	13363 : 0;
	13364 : 0;
	13365 : 1;
	13366 : 1;
	13367 : 1;
	13368 : 0;
	13369 : 1;
	13370 : 0;
	13371 : 1;
	13372 : 1;
	13373 : 0;
	13374 : 1;
	13375 : 1;
	13376 : 0;
	13377 : 1;
	13378 : 1;
	13379 : 0;
	13380 : 1;
	13381 : 1;
	13382 : 1;
	13383 : 1;
	13384 : 1;
	13385 : 1;
	13386 : 1;
	13387 : 0;
	13388 : 0;
	13389 : 0;
	13390 : 0;
	13391 : 1;
	13392 : 1;
	13393 : 0;
	13394 : 0;
	13395 : 1;
	13396 : 0;
	13397 : 1;
	13398 : 1;
	13399 : 1;
	13400 : 0;
	13401 : 1;
	13402 : 0;
	13403 : 1;
	13404 : 1;
	13405 : 0;
	13406 : 1;
	13407 : 1;
	13408 : 1;
	13409 : 1;
	13410 : 1;
	13411 : 1;
	13412 : 1;
	13413 : 1;
	13414 : 1;
	13415 : 1;
	13416 : 1;
	13417 : 1;
	13418 : 1;
	13419 : 1;
	13420 : 1;
	13421 : 1;
	13422 : 1;
	13423 : 1;
	13424 : 1;
	13425 : 1;
	13426 : 1;
	13427 : 1;
	13428 : 1;
	13429 : 1;
	13430 : 1;
	13431 : 1;
	13432 : 1;
	13433 : 1;
	13434 : 1;
	13435 : 1;
	13436 : 1;
	13437 : 1;
	13438 : 1;
	13439 : 1;
	13440 : 1;
	13441 : 1;
	13442 : 1;
	13443 : 1;
	13444 : 1;
	13445 : 1;
	13446 : 1;
	13447 : 1;
	13448 : 1;
	13449 : 1;
	13450 : 1;
	13451 : 1;
	13452 : 1;
	13453 : 1;
	13454 : 1;
	13455 : 1;
	13456 : 1;
	13457 : 1;
	13458 : 1;
	13459 : 1;
	13460 : 1;
	13461 : 1;
	13462 : 1;
	13463 : 1;
	13464 : 1;
	13465 : 1;
	13466 : 1;
	13467 : 1;
	13468 : 1;
	13469 : 1;
	13470 : 1;
	13471 : 1;
	13472 : 1;
	13473 : 0;
	13474 : 0;
	13475 : 0;
	13476 : 0;
	13477 : 1;
	13478 : 1;
	13479 : 1;
	13480 : 0;
	13481 : 1;
	13482 : 0;
	13483 : 0;
	13484 : 0;
	13485 : 0;
	13486 : 0;
	13487 : 1;
	13488 : 0;
	13489 : 1;
	13490 : 1;
	13491 : 1;
	13492 : 1;
	13493 : 1;
	13494 : 0;
	13495 : 1;
	13496 : 0;
	13497 : 1;
	13498 : 1;
	13499 : 1;
	13500 : 0;
	13501 : 0;
	13502 : 1;
	13503 : 0;
	13504 : 0;
	13505 : 1;
	13506 : 1;
	13507 : 1;
	13508 : 1;
	13509 : 0;
	13510 : 1;
	13511 : 1;
	13512 : 1;
	13513 : 0;
	13514 : 1;
	13515 : 1;
	13516 : 1;
	13517 : 0;
	13518 : 1;
	13519 : 0;
	13520 : 1;
	13521 : 1;
	13522 : 1;
	13523 : 0;
	13524 : 0;
	13525 : 0;
	13526 : 0;
	13527 : 1;
	13528 : 0;
	13529 : 0;
	13530 : 1;
	13531 : 0;
	13532 : 0;
	13533 : 1;
	13534 : 1;
	13535 : 1;
	13536 : 1;
	13537 : 0;
	13538 : 0;
	13539 : 1;
	13540 : 1;
	13541 : 1;
	13542 : 1;
	13543 : 1;
	13544 : 0;
	13545 : 1;
	13546 : 1;
	13547 : 1;
	13548 : 0;
	13549 : 1;
	13550 : 1;
	13551 : 1;
	13552 : 0;
	13553 : 0;
	13554 : 1;
	13555 : 1;
	13556 : 1;
	13557 : 0;
	13558 : 1;
	13559 : 1;
	13560 : 1;
	13561 : 0;
	13562 : 1;
	13563 : 0;
	13564 : 1;
	13565 : 1;
	13566 : 0;
	13567 : 1;
	13568 : 1;
	13569 : 0;
	13570 : 1;
	13571 : 1;
	13572 : 1;
	13573 : 1;
	13574 : 1;
	13575 : 1;
	13576 : 1;
	13577 : 1;
	13578 : 0;
	13579 : 0;
	13580 : 1;
	13581 : 1;
	13582 : 1;
	13583 : 0;
	13584 : 1;
	13585 : 1;
	13586 : 1;
	13587 : 0;
	13588 : 1;
	13589 : 1;
	13590 : 1;
	13591 : 0;
	13592 : 1;
	13593 : 1;
	13594 : 1;
	13595 : 0;
	13596 : 1;
	13597 : 0;
	13598 : 1;
	13599 : 1;
	13600 : 1;
	13601 : 0;
	13602 : 0;
	13603 : 0;
	13604 : 0;
	13605 : 1;
	13606 : 1;
	13607 : 1;
	13608 : 0;
	13609 : 1;
	13610 : 0;
	13611 : 1;
	13612 : 1;
	13613 : 0;
	13614 : 1;
	13615 : 1;
	13616 : 0;
	13617 : 1;
	13618 : 1;
	13619 : 0;
	13620 : 1;
	13621 : 1;
	13622 : 1;
	13623 : 1;
	13624 : 1;
	13625 : 1;
	13626 : 1;
	13627 : 0;
	13628 : 0;
	13629 : 0;
	13630 : 0;
	13631 : 0;
	13632 : 0;
	13633 : 0;
	13634 : 0;
	13635 : 1;
	13636 : 0;
	13637 : 1;
	13638 : 1;
	13639 : 1;
	13640 : 0;
	13641 : 1;
	13642 : 0;
	13643 : 1;
	13644 : 1;
	13645 : 0;
	13646 : 1;
	13647 : 1;
	13648 : 1;
	13649 : 1;
	13650 : 1;
	13651 : 1;
	13652 : 1;
	13653 : 1;
	13654 : 1;
	13655 : 1;
	13656 : 1;
	13657 : 1;
	13658 : 1;
	13659 : 1;
	13660 : 1;
	13661 : 1;
	13662 : 1;
	13663 : 1;
	13664 : 1;
	13665 : 1;
	13666 : 1;
	13667 : 1;
	13668 : 1;
	13669 : 1;
	13670 : 1;
	13671 : 1;
	13672 : 1;
	13673 : 1;
	13674 : 1;
	13675 : 1;
	13676 : 1;
	13677 : 1;
	13678 : 1;
	13679 : 1;
	13680 : 1;
	13681 : 1;
	13682 : 1;
	13683 : 1;
	13684 : 1;
	13685 : 1;
	13686 : 1;
	13687 : 1;
	13688 : 1;
	13689 : 1;
	13690 : 1;
	13691 : 1;
	13692 : 1;
	13693 : 1;
	13694 : 1;
	13695 : 1;
	13696 : 1;
	13697 : 1;
	13698 : 1;
	13699 : 1;
	13700 : 1;
	13701 : 1;
	13702 : 1;
	13703 : 1;
	13704 : 1;
	13705 : 1;
	13706 : 1;
	13707 : 1;
	13708 : 1;
	13709 : 0;
	13710 : 1;
	13711 : 1;
	13712 : 1;
	13713 : 0;
	13714 : 0;
	13715 : 0;
	13716 : 0;
	13717 : 1;
	13718 : 1;
	13719 : 1;
	13720 : 0;
	13721 : 1;
	13722 : 0;
	13723 : 1;
	13724 : 1;
	13725 : 1;
	13726 : 1;
	13727 : 1;
	13728 : 0;
	13729 : 1;
	13730 : 1;
	13731 : 1;
	13732 : 0;
	13733 : 1;
	13734 : 0;
	13735 : 1;
	13736 : 0;
	13737 : 1;
	13738 : 1;
	13739 : 0;
	13740 : 0;
	13741 : 0;
	13742 : 1;
	13743 : 0;
	13744 : 0;
	13745 : 1;
	13746 : 1;
	13747 : 1;
	13748 : 1;
	13749 : 0;
	13750 : 1;
	13751 : 1;
	13752 : 1;
	13753 : 0;
	13754 : 1;
	13755 : 1;
	13756 : 1;
	13757 : 0;
	13758 : 1;
	13759 : 0;
	13760 : 1;
	13761 : 1;
	13762 : 0;
	13763 : 0;
	13764 : 0;
	13765 : 0;
	13766 : 0;
	13767 : 1;
	13768 : 0;
	13769 : 0;
	13770 : 1;
	13771 : 0;
	13772 : 1;
	13773 : 0;
	13774 : 1;
	13775 : 1;
	13776 : 1;
	13777 : 1;
	13778 : 1;
	13779 : 0;
	13780 : 1;
	13781 : 1;
	13782 : 1;
	13783 : 1;
	13784 : 0;
	13785 : 1;
	13786 : 1;
	13787 : 1;
	13788 : 0;
	13789 : 1;
	13790 : 1;
	13791 : 1;
	13792 : 0;
	13793 : 0;
	13794 : 1;
	13795 : 1;
	13796 : 1;
	13797 : 0;
	13798 : 1;
	13799 : 1;
	13800 : 1;
	13801 : 0;
	13802 : 1;
	13803 : 0;
	13804 : 1;
	13805 : 1;
	13806 : 0;
	13807 : 1;
	13808 : 1;
	13809 : 0;
	13810 : 1;
	13811 : 1;
	13812 : 1;
	13813 : 1;
	13814 : 1;
	13815 : 1;
	13816 : 1;
	13817 : 1;
	13818 : 0;
	13819 : 0;
	13820 : 1;
	13821 : 1;
	13822 : 1;
	13823 : 0;
	13824 : 1;
	13825 : 1;
	13826 : 1;
	13827 : 0;
	13828 : 1;
	13829 : 1;
	13830 : 1;
	13831 : 0;
	13832 : 1;
	13833 : 1;
	13834 : 1;
	13835 : 0;
	13836 : 1;
	13837 : 0;
	13838 : 1;
	13839 : 1;
	13840 : 1;
	13841 : 0;
	13842 : 0;
	13843 : 0;
	13844 : 0;
	13845 : 1;
	13846 : 1;
	13847 : 1;
	13848 : 0;
	13849 : 1;
	13850 : 0;
	13851 : 1;
	13852 : 1;
	13853 : 0;
	13854 : 1;
	13855 : 1;
	13856 : 0;
	13857 : 1;
	13858 : 1;
	13859 : 0;
	13860 : 1;
	13861 : 1;
	13862 : 1;
	13863 : 0;
	13864 : 1;
	13865 : 1;
	13866 : 1;
	13867 : 0;
	13868 : 0;
	13869 : 0;
	13870 : 0;
	13871 : 1;
	13872 : 1;
	13873 : 1;
	13874 : 1;
	13875 : 1;
	13876 : 0;
	13877 : 1;
	13878 : 1;
	13879 : 1;
	13880 : 0;
	13881 : 1;
	13882 : 0;
	13883 : 1;
	13884 : 1;
	13885 : 0;
	13886 : 1;
	13887 : 0;
	13888 : 0;
	13889 : 1;
	13890 : 1;
	13891 : 1;
	13892 : 1;
	13893 : 1;
	13894 : 1;
	13895 : 1;
	13896 : 1;
	13897 : 1;
	13898 : 1;
	13899 : 1;
	13900 : 1;
	13901 : 1;
	13902 : 1;
	13903 : 1;
	13904 : 1;
	13905 : 1;
	13906 : 1;
	13907 : 1;
	13908 : 1;
	13909 : 1;
	13910 : 1;
	13911 : 1;
	13912 : 1;
	13913 : 1;
	13914 : 1;
	13915 : 1;
	13916 : 1;
	13917 : 1;
	13918 : 1;
	13919 : 1;
	13920 : 1;
	13921 : 1;
	13922 : 1;
	13923 : 1;
	13924 : 1;
	13925 : 1;
	13926 : 1;
	13927 : 1;
	13928 : 1;
	13929 : 1;
	13930 : 1;
	13931 : 1;
	13932 : 1;
	13933 : 1;
	13934 : 1;
	13935 : 1;
	13936 : 1;
	13937 : 1;
	13938 : 1;
	13939 : 1;
	13940 : 1;
	13941 : 1;
	13942 : 1;
	13943 : 1;
	13944 : 1;
	13945 : 1;
	13946 : 1;
	13947 : 1;
	13948 : 1;
	13949 : 1;
	13950 : 0;
	13951 : 0;
	13952 : 0;
	13953 : 0;
	13954 : 1;
	13955 : 0;
	13956 : 0;
	13957 : 0;
	13958 : 0;
	13959 : 0;
	13960 : 1;
	13961 : 1;
	13962 : 1;
	13963 : 0;
	13964 : 0;
	13965 : 0;
	13966 : 0;
	13967 : 1;
	13968 : 1;
	13969 : 0;
	13970 : 0;
	13971 : 0;
	13972 : 1;
	13973 : 1;
	13974 : 0;
	13975 : 1;
	13976 : 1;
	13977 : 0;
	13978 : 0;
	13979 : 0;
	13980 : 0;
	13981 : 0;
	13982 : 1;
	13983 : 0;
	13984 : 0;
	13985 : 1;
	13986 : 1;
	13987 : 1;
	13988 : 1;
	13989 : 0;
	13990 : 0;
	13991 : 0;
	13992 : 1;
	13993 : 0;
	13994 : 1;
	13995 : 1;
	13996 : 1;
	13997 : 0;
	13998 : 1;
	13999 : 1;
	14000 : 0;
	14001 : 0;
	14002 : 0;
	14003 : 0;
	14004 : 0;
	14005 : 0;
	14006 : 0;
	14007 : 1;
	14008 : 0;
	14009 : 0;
	14010 : 1;
	14011 : 0;
	14012 : 1;
	14013 : 1;
	14014 : 0;
	14015 : 1;
	14016 : 0;
	14017 : 0;
	14018 : 0;
	14019 : 0;
	14020 : 1;
	14021 : 1;
	14022 : 1;
	14023 : 1;
	14024 : 0;
	14025 : 0;
	14026 : 0;
	14027 : 0;
	14028 : 1;
	14029 : 0;
	14030 : 0;
	14031 : 0;
	14032 : 0;
	14033 : 1;
	14034 : 1;
	14035 : 1;
	14036 : 1;
	14037 : 1;
	14038 : 0;
	14039 : 0;
	14040 : 0;
	14041 : 1;
	14042 : 1;
	14043 : 1;
	14044 : 0;
	14045 : 0;
	14046 : 1;
	14047 : 0;
	14048 : 1;
	14049 : 0;
	14050 : 1;
	14051 : 1;
	14052 : 1;
	14053 : 1;
	14054 : 1;
	14055 : 1;
	14056 : 1;
	14057 : 1;
	14058 : 0;
	14059 : 0;
	14060 : 1;
	14061 : 1;
	14062 : 1;
	14063 : 0;
	14064 : 1;
	14065 : 1;
	14066 : 1;
	14067 : 0;
	14068 : 1;
	14069 : 1;
	14070 : 1;
	14071 : 0;
	14072 : 0;
	14073 : 0;
	14074 : 0;
	14075 : 1;
	14076 : 1;
	14077 : 1;
	14078 : 0;
	14079 : 0;
	14080 : 0;
	14081 : 0;
	14082 : 1;
	14083 : 0;
	14084 : 0;
	14085 : 1;
	14086 : 1;
	14087 : 1;
	14088 : 0;
	14089 : 1;
	14090 : 1;
	14091 : 0;
	14092 : 0;
	14093 : 1;
	14094 : 0;
	14095 : 1;
	14096 : 0;
	14097 : 1;
	14098 : 1;
	14099 : 0;
	14100 : 1;
	14101 : 1;
	14102 : 1;
	14103 : 1;
	14104 : 0;
	14105 : 0;
	14106 : 0;
	14107 : 0;
	14108 : 1;
	14109 : 1;
	14110 : 0;
	14111 : 0;
	14112 : 0;
	14113 : 0;
	14114 : 0;
	14115 : 1;
	14116 : 1;
	14117 : 0;
	14118 : 0;
	14119 : 0;
	14120 : 1;
	14121 : 1;
	14122 : 0;
	14123 : 1;
	14124 : 1;
	14125 : 0;
	14126 : 1;
	14127 : 0;
	14128 : 0;
	14129 : 1;
	14130 : 1;
	14131 : 1;
	14132 : 1;
	14133 : 1;
	14134 : 1;
	14135 : 1;
	14136 : 1;
	14137 : 1;
	14138 : 1;
	14139 : 1;
	14140 : 1;
	14141 : 1;
	14142 : 1;
	14143 : 1;
	14144 : 1;
	14145 : 1;
	14146 : 1;
	14147 : 1;
	14148 : 1;
	14149 : 1;
	14150 : 1;
	14151 : 1;
	14152 : 1;
	14153 : 1;
	14154 : 1;
	14155 : 1;
	14156 : 1;
	14157 : 1;
	14158 : 1;
	14159 : 1;
	14160 : 1;
	14161 : 1;
	14162 : 1;
	14163 : 1;
	14164 : 1;
	14165 : 1;
	14166 : 1;
	14167 : 1;
	14168 : 1;
	14169 : 1;
	14170 : 1;
	14171 : 1;
	14172 : 1;
	14173 : 1;
	14174 : 1;
	14175 : 1;
	14176 : 1;
	14177 : 1;
	14178 : 1;
	14179 : 1;
	14180 : 1;
	14181 : 1;
	14182 : 1;
	14183 : 1;
	14184 : 1;
	14185 : 1;
	14186 : 1;
	14187 : 1;
	14188 : 1;
	14189 : 1;
	14190 : 1;
	14191 : 1;
	14192 : 1;
	14193 : 1;
	14194 : 1;
	14195 : 0;
	14196 : 0;
	14197 : 1;
	14198 : 1;
	14199 : 1;
	14200 : 1;
	14201 : 1;
	14202 : 1;
	14203 : 1;
	14204 : 1;
	14205 : 1;
	14206 : 1;
	14207 : 1;
	14208 : 1;
	14209 : 1;
	14210 : 1;
	14211 : 1;
	14212 : 1;
	14213 : 1;
	14214 : 1;
	14215 : 1;
	14216 : 1;
	14217 : 1;
	14218 : 1;
	14219 : 1;
	14220 : 1;
	14221 : 1;
	14222 : 1;
	14223 : 1;
	14224 : 1;
	14225 : 1;
	14226 : 1;
	14227 : 1;
	14228 : 1;
	14229 : 1;
	14230 : 1;
	14231 : 1;
	14232 : 1;
	14233 : 1;
	14234 : 1;
	14235 : 1;
	14236 : 1;
	14237 : 1;
	14238 : 1;
	14239 : 1;
	14240 : 1;
	14241 : 1;
	14242 : 1;
	14243 : 1;
	14244 : 1;
	14245 : 1;
	14246 : 1;
	14247 : 1;
	14248 : 1;
	14249 : 1;
	14250 : 1;
	14251 : 1;
	14252 : 1;
	14253 : 1;
	14254 : 1;
	14255 : 1;
	14256 : 1;
	14257 : 1;
	14258 : 1;
	14259 : 1;
	14260 : 1;
	14261 : 1;
	14262 : 1;
	14263 : 1;
	14264 : 1;
	14265 : 1;
	14266 : 1;
	14267 : 1;
	14268 : 1;
	14269 : 1;
	14270 : 1;
	14271 : 1;
	14272 : 1;
	14273 : 1;
	14274 : 1;
	14275 : 1;
	14276 : 1;
	14277 : 1;
	14278 : 1;
	14279 : 1;
	14280 : 1;
	14281 : 1;
	14282 : 1;
	14283 : 1;
	14284 : 1;
	14285 : 1;
	14286 : 1;
	14287 : 1;
	14288 : 1;
	14289 : 1;
	14290 : 1;
	14291 : 1;
	14292 : 1;
	14293 : 1;
	14294 : 1;
	14295 : 1;
	14296 : 1;
	14297 : 1;
	14298 : 1;
	14299 : 1;
	14300 : 1;
	14301 : 1;
	14302 : 1;
	14303 : 1;
	14304 : 1;
	14305 : 1;
	14306 : 1;
	14307 : 1;
	14308 : 1;
	14309 : 1;
	14310 : 1;
	14311 : 1;
	14312 : 1;
	14313 : 1;
	14314 : 1;
	14315 : 1;
	14316 : 1;
	14317 : 1;
	14318 : 1;
	14319 : 1;
	14320 : 1;
	14321 : 1;
	14322 : 1;
	14323 : 1;
	14324 : 1;
	14325 : 1;
	14326 : 1;
	14327 : 1;
	14328 : 1;
	14329 : 1;
	14330 : 1;
	14331 : 1;
	14332 : 1;
	14333 : 1;
	14334 : 1;
	14335 : 1;
	14336 : 1;
	14337 : 1;
	14338 : 1;
	14339 : 1;
	14340 : 1;
	14341 : 1;
	14342 : 1;
	14343 : 1;
	14344 : 1;
	14345 : 1;
	14346 : 1;
	14347 : 1;
	14348 : 1;
	14349 : 1;
	14350 : 1;
	14351 : 1;
	14352 : 1;
	14353 : 1;
	14354 : 1;
	14355 : 1;
	14356 : 1;
	14357 : 1;
	14358 : 1;
	14359 : 1;
	14360 : 1;
	14361 : 1;
	14362 : 1;
	14363 : 1;
	14364 : 1;
	14365 : 1;
	14366 : 1;
	14367 : 1;
	14368 : 0;
	14369 : 1;
	14370 : 1;
	14371 : 1;
	14372 : 1;
	14373 : 1;
	14374 : 1;
	14375 : 1;
	14376 : 1;
	14377 : 1;
	14378 : 1;
	14379 : 1;
	14380 : 1;
	14381 : 1;
	14382 : 1;
	14383 : 1;
	14384 : 1;
	14385 : 1;
	14386 : 1;
	14387 : 1;
	14388 : 1;
	14389 : 1;
	14390 : 1;
	14391 : 1;
	14392 : 1;
	14393 : 1;
	14394 : 1;
	14395 : 1;
	14396 : 1;
	14397 : 1;
	14398 : 1;
	14399 : 1;
	14400 : 1;
	14401 : 1;
	14402 : 1;
	14403 : 1;
	14404 : 1;
	14405 : 1;
	14406 : 1;
	14407 : 1;
	14408 : 1;
	14409 : 1;
	14410 : 1;
	14411 : 1;
	14412 : 1;
	14413 : 1;
	14414 : 1;
	14415 : 1;
	14416 : 1;
	14417 : 1;
	14418 : 1;
	14419 : 1;
	14420 : 1;
	14421 : 1;
	14422 : 1;
	14423 : 1;
	14424 : 1;
	14425 : 1;
	14426 : 1;
	14427 : 1;
	14428 : 1;
	14429 : 1;
	14430 : 1;
	14431 : 1;
	14432 : 1;
	14433 : 1;
	14434 : 1;
	14435 : 0;
	14436 : 0;
	14437 : 1;
	14438 : 1;
	14439 : 1;
	14440 : 1;
	14441 : 1;
	14442 : 1;
	14443 : 1;
	14444 : 1;
	14445 : 1;
	14446 : 1;
	14447 : 1;
	14448 : 1;
	14449 : 1;
	14450 : 1;
	14451 : 1;
	14452 : 1;
	14453 : 1;
	14454 : 1;
	14455 : 1;
	14456 : 1;
	14457 : 1;
	14458 : 1;
	14459 : 1;
	14460 : 1;
	14461 : 1;
	14462 : 1;
	14463 : 1;
	14464 : 1;
	14465 : 1;
	14466 : 1;
	14467 : 1;
	14468 : 1;
	14469 : 1;
	14470 : 1;
	14471 : 1;
	14472 : 1;
	14473 : 1;
	14474 : 1;
	14475 : 1;
	14476 : 1;
	14477 : 1;
	14478 : 1;
	14479 : 1;
	14480 : 1;
	14481 : 1;
	14482 : 1;
	14483 : 1;
	14484 : 1;
	14485 : 1;
	14486 : 1;
	14487 : 1;
	14488 : 1;
	14489 : 1;
	14490 : 1;
	14491 : 1;
	14492 : 1;
	14493 : 1;
	14494 : 1;
	14495 : 1;
	14496 : 1;
	14497 : 1;
	14498 : 1;
	14499 : 1;
	14500 : 1;
	14501 : 1;
	14502 : 1;
	14503 : 1;
	14504 : 1;
	14505 : 1;
	14506 : 1;
	14507 : 1;
	14508 : 1;
	14509 : 1;
	14510 : 1;
	14511 : 1;
	14512 : 1;
	14513 : 1;
	14514 : 1;
	14515 : 1;
	14516 : 1;
	14517 : 1;
	14518 : 1;
	14519 : 1;
	14520 : 1;
	14521 : 1;
	14522 : 1;
	14523 : 1;
	14524 : 1;
	14525 : 1;
	14526 : 1;
	14527 : 1;
	14528 : 1;
	14529 : 1;
	14530 : 1;
	14531 : 1;
	14532 : 1;
	14533 : 1;
	14534 : 1;
	14535 : 1;
	14536 : 1;
	14537 : 1;
	14538 : 1;
	14539 : 1;
	14540 : 1;
	14541 : 1;
	14542 : 1;
	14543 : 1;
	14544 : 1;
	14545 : 1;
	14546 : 1;
	14547 : 1;
	14548 : 1;
	14549 : 1;
	14550 : 1;
	14551 : 1;
	14552 : 1;
	14553 : 1;
	14554 : 1;
	14555 : 1;
	14556 : 1;
	14557 : 1;
	14558 : 1;
	14559 : 1;
	14560 : 1;
	14561 : 1;
	14562 : 1;
	14563 : 1;
	14564 : 1;
	14565 : 1;
	14566 : 1;
	14567 : 1;
	14568 : 1;
	14569 : 1;
	14570 : 1;
	14571 : 1;
	14572 : 1;
	14573 : 1;
	14574 : 1;
	14575 : 1;
	14576 : 1;
	14577 : 1;
	14578 : 1;
	14579 : 1;
	14580 : 1;
	14581 : 1;
	14582 : 1;
	14583 : 1;
	14584 : 1;
	14585 : 1;
	14586 : 1;
	14587 : 1;
	14588 : 1;
	14589 : 1;
	14590 : 1;
	14591 : 1;
	14592 : 1;
	14593 : 1;
	14594 : 1;
	14595 : 1;
	14596 : 1;
	14597 : 1;
	14598 : 1;
	14599 : 1;
	14600 : 1;
	14601 : 1;
	14602 : 1;
	14603 : 1;
	14604 : 1;
	14605 : 1;
	14606 : 1;
	14607 : 0;
	14608 : 1;
	14609 : 1;
	14610 : 1;
	14611 : 1;
	14612 : 1;
	14613 : 1;
	14614 : 1;
	14615 : 1;
	14616 : 1;
	14617 : 1;
	14618 : 1;
	14619 : 1;
	14620 : 1;
	14621 : 1;
	14622 : 1;
	14623 : 1;
	14624 : 1;
	14625 : 1;
	14626 : 1;
	14627 : 1;
	14628 : 1;
	14629 : 1;
	14630 : 1;
	14631 : 1;
	14632 : 1;
	14633 : 1;
	14634 : 1;
	14635 : 1;
	14636 : 1;
	14637 : 1;
	14638 : 1;
	14639 : 1;
	14640 : 1;
	14641 : 1;
	14642 : 1;
	14643 : 1;
	14644 : 1;
	14645 : 1;
	14646 : 1;
	14647 : 1;
	14648 : 1;
	14649 : 1;
	14650 : 1;
	14651 : 1;
	14652 : 1;
	14653 : 1;
	14654 : 1;
	14655 : 1;
	14656 : 1;
	14657 : 1;
	14658 : 1;
	14659 : 1;
	14660 : 1;
	14661 : 1;
	14662 : 1;
	14663 : 1;
	14664 : 1;
	14665 : 1;
	14666 : 1;
	14667 : 1;
	14668 : 1;
	14669 : 1;
	14670 : 1;
	14671 : 1;
	14672 : 1;
	14673 : 1;
	14674 : 1;
	14675 : 1;
	14676 : 1;
	14677 : 1;
	14678 : 1;
	14679 : 1;
	14680 : 1;
	14681 : 1;
	14682 : 1;
	14683 : 1;
	14684 : 1;
	14685 : 1;
	14686 : 1;
	14687 : 1;
	14688 : 1;
	14689 : 1;
	14690 : 1;
	14691 : 1;
	14692 : 1;
	14693 : 1;
	14694 : 1;
	14695 : 1;
	14696 : 1;
	14697 : 1;
	14698 : 1;
	14699 : 1;
	14700 : 1;
	14701 : 1;
	14702 : 1;
	14703 : 1;
	14704 : 1;
	14705 : 1;
	14706 : 1;
	14707 : 1;
	14708 : 1;
	14709 : 1;
	14710 : 1;
	14711 : 1;
	14712 : 1;
	14713 : 1;
	14714 : 1;
	14715 : 1;
	14716 : 1;
	14717 : 1;
	14718 : 1;
	14719 : 1;
	14720 : 1;
	14721 : 1;
	14722 : 1;
	14723 : 1;
	14724 : 1;
	14725 : 1;
	14726 : 1;
	14727 : 1;
	14728 : 1;
	14729 : 1;
	14730 : 1;
	14731 : 1;
	14732 : 1;
	14733 : 1;
	14734 : 1;
	14735 : 1;
	14736 : 1;
	14737 : 1;
	14738 : 1;
	14739 : 1;
	14740 : 1;
	14741 : 1;
	14742 : 1;
	14743 : 1;
	14744 : 1;
	14745 : 1;
	14746 : 1;
	14747 : 1;
	14748 : 1;
	14749 : 1;
	14750 : 1;
	14751 : 1;
	14752 : 1;
	14753 : 1;
	14754 : 1;
	14755 : 1;
	14756 : 1;
	14757 : 1;
	14758 : 1;
	14759 : 1;
	14760 : 1;
	14761 : 1;
	14762 : 1;
	14763 : 1;
	14764 : 1;
	14765 : 1;
	14766 : 1;
	14767 : 1;
	14768 : 1;
	14769 : 1;
	14770 : 1;
	14771 : 1;
	14772 : 1;
	14773 : 1;
	14774 : 1;
	14775 : 1;
	14776 : 1;
	14777 : 1;
	14778 : 1;
	14779 : 1;
	14780 : 1;
	14781 : 1;
	14782 : 1;
	14783 : 1;
	14784 : 1;
	14785 : 1;
	14786 : 1;
	14787 : 1;
	14788 : 1;
	14789 : 1;
	14790 : 1;
	14791 : 1;
	14792 : 1;
	14793 : 1;
	14794 : 1;
	14795 : 1;
	14796 : 1;
	14797 : 1;
	14798 : 1;
	14799 : 1;
	14800 : 1;
	14801 : 1;
	14802 : 1;
	14803 : 1;
	14804 : 1;
	14805 : 1;
	14806 : 1;
	14807 : 1;
	14808 : 1;
	14809 : 1;
	14810 : 1;
	14811 : 1;
	14812 : 1;
	14813 : 1;
	14814 : 1;
	14815 : 1;
	14816 : 1;
	14817 : 1;
	14818 : 1;
	14819 : 1;
	14820 : 1;
	14821 : 1;
	14822 : 1;
	14823 : 1;
	14824 : 1;
	14825 : 1;
	14826 : 1;
	14827 : 1;
	14828 : 1;
	14829 : 1;
	14830 : 1;
	14831 : 1;
	14832 : 1;
	14833 : 1;
	14834 : 1;
	14835 : 1;
	14836 : 1;
	14837 : 1;
	14838 : 1;
	14839 : 1;
	14840 : 1;
	14841 : 1;
	14842 : 1;
	14843 : 1;
	14844 : 1;
	14845 : 1;
	14846 : 1;
	14847 : 1;
	14848 : 1;
	14849 : 1;
	14850 : 1;
	14851 : 1;
	14852 : 1;
	14853 : 1;
	14854 : 1;
	14855 : 1;
	14856 : 1;
	14857 : 1;
	14858 : 1;
	14859 : 1;
	14860 : 1;
	14861 : 1;
	14862 : 1;
	14863 : 1;
	14864 : 1;
	14865 : 1;
	14866 : 1;
	14867 : 1;
	14868 : 1;
	14869 : 1;
	14870 : 1;
	14871 : 1;
	14872 : 1;
	14873 : 1;
	14874 : 1;
	14875 : 1;
	14876 : 1;
	14877 : 1;
	14878 : 1;
	14879 : 1;
	14880 : 1;
	14881 : 1;
	14882 : 1;
	14883 : 1;
	14884 : 1;
	14885 : 1;
	14886 : 1;
	14887 : 1;
	14888 : 1;
	14889 : 1;
	14890 : 1;
	14891 : 1;
	14892 : 1;
	14893 : 1;
	14894 : 1;
	14895 : 1;
	14896 : 1;
	14897 : 1;
	14898 : 1;
	14899 : 1;
	14900 : 1;
	14901 : 1;
	14902 : 1;
	14903 : 1;
	14904 : 1;
	14905 : 1;
	14906 : 1;
	14907 : 1;
	14908 : 1;
	14909 : 1;
	14910 : 1;
	14911 : 1;
	14912 : 1;
	14913 : 1;
	14914 : 1;
	14915 : 1;
	14916 : 1;
	14917 : 1;
	14918 : 1;
	14919 : 1;
	14920 : 1;
	14921 : 1;
	14922 : 1;
	14923 : 1;
	14924 : 1;
	14925 : 1;
	14926 : 1;
	14927 : 1;
	14928 : 1;
	14929 : 1;
	14930 : 1;
	14931 : 1;
	14932 : 1;
	14933 : 1;
	14934 : 1;
	14935 : 1;
	14936 : 1;
	14937 : 1;
	14938 : 1;
	14939 : 1;
	14940 : 1;
	14941 : 1;
	14942 : 1;
	14943 : 1;
	14944 : 1;
	14945 : 1;
	14946 : 1;
	14947 : 1;
	14948 : 1;
	14949 : 1;
	14950 : 1;
	14951 : 1;
	14952 : 1;
	14953 : 1;
	14954 : 1;
	14955 : 1;
	14956 : 1;
	14957 : 1;
	14958 : 1;
	14959 : 1;
	14960 : 1;
	14961 : 1;
	14962 : 1;
	14963 : 1;
	14964 : 1;
	14965 : 1;
	14966 : 1;
	14967 : 1;
	14968 : 1;
	14969 : 1;
	14970 : 1;
	14971 : 1;
	14972 : 1;
	14973 : 1;
	14974 : 1;
	14975 : 1;
	14976 : 1;
	14977 : 1;
	14978 : 1;
	14979 : 1;
	14980 : 1;
	14981 : 1;
	14982 : 1;
	14983 : 1;
	14984 : 1;
	14985 : 1;
	14986 : 1;
	14987 : 1;
	14988 : 1;
	14989 : 1;
	14990 : 1;
	14991 : 1;
	14992 : 1;
	14993 : 1;
	14994 : 1;
	14995 : 1;
	14996 : 1;
	14997 : 1;
	14998 : 1;
	14999 : 1;
	15000 : 1;
	15001 : 1;
	15002 : 1;
	15003 : 1;
	15004 : 1;
	15005 : 1;
	15006 : 1;
	15007 : 1;
	15008 : 1;
	15009 : 1;
	15010 : 1;
	15011 : 1;
	15012 : 1;
	15013 : 1;
	15014 : 1;
	15015 : 1;
	15016 : 1;
	15017 : 1;
	15018 : 1;
	15019 : 1;
	15020 : 1;
	15021 : 1;
	15022 : 1;
	15023 : 1;
	15024 : 1;
	15025 : 1;
	15026 : 1;
	15027 : 1;
	15028 : 1;
	15029 : 1;
	15030 : 1;
	15031 : 1;
	15032 : 1;
	15033 : 1;
	15034 : 1;
	15035 : 1;
	15036 : 1;
	15037 : 1;
	15038 : 1;
	15039 : 1;
	15040 : 1;
	15041 : 1;
	15042 : 1;
	15043 : 1;
	15044 : 1;
	15045 : 1;
	15046 : 1;
	15047 : 1;
	15048 : 1;
	15049 : 1;
	15050 : 1;
	15051 : 1;
	15052 : 1;
	15053 : 1;
	15054 : 1;
	15055 : 1;
	15056 : 1;
	15057 : 1;
	15058 : 1;
	15059 : 1;
	15060 : 1;
	15061 : 1;
	15062 : 1;
	15063 : 1;
	15064 : 1;
	15065 : 1;
	15066 : 1;
	15067 : 1;
	15068 : 1;
	15069 : 1;
	15070 : 1;
	15071 : 1;
	15072 : 1;
	15073 : 1;
	15074 : 1;
	15075 : 1;
	15076 : 1;
	15077 : 1;
	15078 : 1;
	15079 : 1;
	15080 : 1;
	15081 : 1;
	15082 : 1;
	15083 : 1;
	15084 : 1;
	15085 : 1;
	15086 : 1;
	15087 : 1;
	15088 : 1;
	15089 : 1;
	15090 : 1;
	15091 : 1;
	15092 : 1;
	15093 : 1;
	15094 : 1;
	15095 : 1;
	15096 : 1;
	15097 : 1;
	15098 : 1;
	15099 : 1;
	15100 : 1;
	15101 : 1;
	15102 : 1;
	15103 : 1;
	15104 : 1;
	15105 : 1;
	15106 : 1;
	15107 : 1;
	15108 : 1;
	15109 : 1;
	15110 : 1;
	15111 : 1;
	15112 : 1;
	15113 : 1;
	15114 : 1;
	15115 : 1;
	15116 : 1;
	15117 : 1;
	15118 : 1;
	15119 : 1;
	15120 : 1;
	15121 : 1;
	15122 : 1;
	15123 : 1;
	15124 : 1;
	15125 : 1;
	15126 : 1;
	15127 : 1;
	15128 : 1;
	15129 : 1;
	15130 : 1;
	15131 : 1;
	15132 : 1;
	15133 : 1;
	15134 : 1;
	15135 : 1;
	15136 : 1;
	15137 : 1;
	15138 : 1;
	15139 : 1;
	15140 : 1;
	15141 : 1;
	15142 : 1;
	15143 : 1;
	15144 : 1;
	15145 : 1;
	15146 : 1;
	15147 : 1;
	15148 : 1;
	15149 : 1;
	15150 : 1;
	15151 : 1;
	15152 : 1;
	15153 : 1;
	15154 : 1;
	15155 : 1;
	15156 : 1;
	15157 : 1;
	15158 : 1;
	15159 : 1;
	15160 : 1;
	15161 : 1;
	15162 : 1;
	15163 : 1;
	15164 : 1;
	15165 : 1;
	15166 : 1;
	15167 : 1;
	15168 : 1;
	15169 : 1;
	15170 : 1;
	15171 : 1;
	15172 : 1;
	15173 : 1;
	15174 : 1;
	15175 : 1;
	15176 : 1;
	15177 : 1;
	15178 : 1;
	15179 : 1;
	15180 : 1;
	15181 : 1;
	15182 : 1;
	15183 : 1;
	15184 : 1;
	15185 : 1;
	15186 : 1;
	15187 : 1;
	15188 : 1;
	15189 : 1;
	15190 : 1;
	15191 : 1;
	15192 : 1;
	15193 : 1;
	15194 : 1;
	15195 : 1;
	15196 : 1;
	15197 : 1;
	15198 : 1;
	15199 : 1;
	15200 : 1;
	15201 : 1;
	15202 : 1;
	15203 : 1;
	15204 : 1;
	15205 : 1;
	15206 : 1;
	15207 : 1;
	15208 : 1;
	15209 : 1;
	15210 : 1;
	15211 : 1;
	15212 : 1;
	15213 : 1;
	15214 : 1;
	15215 : 1;
	15216 : 1;
	15217 : 1;
	15218 : 1;
	15219 : 1;
	15220 : 1;
	15221 : 1;
	15222 : 1;
	15223 : 1;
	15224 : 1;
	15225 : 1;
	15226 : 1;
	15227 : 1;
	15228 : 1;
	15229 : 1;
	15230 : 1;
	15231 : 1;
	15232 : 1;
	15233 : 1;
	15234 : 1;
	15235 : 1;
	15236 : 1;
	15237 : 1;
	15238 : 1;
	15239 : 1;
	15240 : 1;
	15241 : 1;
	15242 : 1;
	15243 : 1;
	15244 : 1;
	15245 : 1;
	15246 : 1;
	15247 : 1;
	15248 : 1;
	15249 : 1;
	15250 : 1;
	15251 : 1;
	15252 : 1;
	15253 : 1;
	15254 : 1;
	15255 : 1;
	15256 : 1;
	15257 : 1;
	15258 : 1;
	15259 : 1;
	15260 : 1;
	15261 : 1;
	15262 : 1;
	15263 : 1;
	15264 : 1;
	15265 : 1;
	15266 : 1;
	15267 : 1;
	15268 : 1;
	15269 : 1;
	15270 : 1;
	15271 : 1;
	15272 : 1;
	15273 : 1;
	15274 : 1;
	15275 : 1;
	15276 : 1;
	15277 : 1;
	15278 : 1;
	15279 : 1;
	15280 : 1;
	15281 : 1;
	15282 : 1;
	15283 : 1;
	15284 : 1;
	15285 : 1;
	15286 : 1;
	15287 : 1;
	15288 : 1;
	15289 : 1;
	15290 : 1;
	15291 : 1;
	15292 : 1;
	15293 : 1;
	15294 : 1;
	15295 : 1;
	15296 : 1;
	15297 : 1;
	15298 : 1;
	15299 : 1;
	15300 : 1;
	15301 : 1;
	15302 : 1;
	15303 : 1;
	15304 : 1;
	15305 : 1;
	15306 : 1;
	15307 : 1;
	15308 : 1;
	15309 : 1;
	15310 : 1;
	15311 : 1;
	15312 : 1;
	15313 : 1;
	15314 : 1;
	15315 : 1;
	15316 : 1;
	15317 : 1;
	15318 : 1;
	15319 : 1;
	15320 : 1;
	15321 : 1;
	15322 : 1;
	15323 : 1;
	15324 : 1;
	15325 : 1;
	15326 : 1;
	15327 : 1;
	15328 : 1;
	15329 : 1;
	15330 : 1;
	15331 : 1;
	15332 : 1;
	15333 : 1;
	15334 : 1;
	15335 : 1;
	15336 : 1;
	15337 : 1;
	15338 : 1;
	15339 : 1;
	15340 : 1;
	15341 : 1;
	15342 : 1;
	15343 : 1;
	15344 : 1;
	15345 : 1;
	15346 : 1;
	15347 : 1;
	15348 : 1;
	15349 : 1;
	15350 : 1;
	15351 : 1;
	15352 : 1;
	15353 : 1;
	15354 : 1;
	15355 : 1;
	15356 : 1;
	15357 : 1;
	15358 : 1;
	15359 : 1;
	15360 : 1;
	15361 : 1;
	15362 : 1;
	15363 : 1;
	15364 : 1;
	15365 : 1;
	15366 : 1;
	15367 : 1;
	15368 : 1;
	15369 : 1;
	15370 : 1;
	15371 : 1;
	15372 : 1;
	15373 : 1;
	15374 : 1;
	15375 : 1;
	15376 : 1;
	15377 : 1;
	15378 : 1;
	15379 : 1;
	15380 : 1;
	15381 : 1;
	15382 : 1;
	15383 : 1;
	15384 : 1;
	15385 : 1;
	15386 : 1;
	15387 : 1;
	15388 : 1;
	15389 : 1;
	15390 : 1;
	15391 : 1;
	15392 : 1;
	15393 : 1;
	15394 : 1;
	15395 : 1;
	15396 : 1;
	15397 : 1;
	15398 : 1;
	15399 : 1;
	15400 : 1;
	15401 : 1;
	15402 : 1;
	15403 : 1;
	15404 : 1;
	15405 : 1;
	15406 : 1;
	15407 : 1;
	15408 : 1;
	15409 : 1;
	15410 : 1;
	15411 : 1;
	15412 : 1;
	15413 : 1;
	15414 : 1;
	15415 : 1;
	15416 : 1;
	15417 : 1;
	15418 : 1;
	15419 : 1;
	15420 : 1;
	15421 : 1;
	15422 : 1;
	15423 : 1;
	15424 : 1;
	15425 : 1;
	15426 : 1;
	15427 : 1;
	15428 : 1;
	15429 : 1;
	15430 : 1;
	15431 : 1;
	15432 : 1;
	15433 : 1;
	15434 : 1;
	15435 : 1;
	15436 : 1;
	15437 : 1;
	15438 : 1;
	15439 : 1;
	15440 : 1;
	15441 : 1;
	15442 : 1;
	15443 : 1;
	15444 : 1;
	15445 : 1;
	15446 : 1;
	15447 : 1;
	15448 : 1;
	15449 : 1;
	15450 : 1;
	15451 : 1;
	15452 : 1;
	15453 : 1;
	15454 : 1;
	15455 : 1;
	15456 : 1;
	15457 : 1;
	15458 : 1;
	15459 : 1;
	15460 : 1;
	15461 : 1;
	15462 : 1;
	15463 : 1;
	15464 : 1;
	15465 : 1;
	15466 : 1;
	15467 : 1;
	15468 : 1;
	15469 : 1;
	15470 : 1;
	15471 : 1;
	15472 : 1;
	15473 : 1;
	15474 : 1;
	15475 : 1;
	15476 : 1;
	15477 : 1;
	15478 : 1;
	15479 : 1;
	15480 : 1;
	15481 : 1;
	15482 : 1;
	15483 : 1;
	15484 : 1;
	15485 : 1;
	15486 : 1;
	15487 : 1;
	15488 : 1;
	15489 : 1;
	15490 : 1;
	15491 : 1;
	15492 : 1;
	15493 : 1;
	15494 : 1;
	15495 : 1;
	15496 : 1;
	15497 : 1;
	15498 : 1;
	15499 : 1;
	15500 : 1;
	15501 : 1;
	15502 : 1;
	15503 : 1;
	15504 : 1;
	15505 : 1;
	15506 : 1;
	15507 : 1;
	15508 : 1;
	15509 : 1;
	15510 : 1;
	15511 : 1;
	15512 : 1;
	15513 : 1;
	15514 : 1;
	15515 : 1;
	15516 : 1;
	15517 : 1;
	15518 : 1;
	15519 : 1;
	15520 : 1;
	15521 : 1;
	15522 : 1;
	15523 : 1;
	15524 : 1;
	15525 : 1;
	15526 : 1;
	15527 : 1;
	15528 : 1;
	15529 : 1;
	15530 : 1;
	15531 : 1;
	15532 : 1;
	15533 : 1;
	15534 : 1;
	15535 : 1;
	15536 : 1;
	15537 : 1;
	15538 : 1;
	15539 : 1;
	15540 : 1;
	15541 : 1;
	15542 : 1;
	15543 : 1;
	15544 : 1;
	15545 : 1;
	15546 : 1;
	15547 : 1;
	15548 : 1;
	15549 : 1;
	15550 : 1;
	15551 : 1;
	15552 : 1;
	15553 : 1;
	15554 : 1;
	15555 : 1;
	15556 : 1;
	15557 : 1;
	15558 : 1;
	15559 : 1;
	15560 : 1;
	15561 : 1;
	15562 : 1;
	15563 : 1;
	15564 : 1;
	15565 : 1;
	15566 : 1;
	15567 : 1;
	15568 : 1;
	15569 : 1;
	15570 : 1;
	15571 : 1;
	15572 : 1;
	15573 : 1;
	15574 : 1;
	15575 : 1;
	15576 : 1;
	15577 : 1;
	15578 : 1;
	15579 : 1;
	15580 : 1;
	15581 : 1;
	15582 : 1;
	15583 : 1;
	15584 : 1;
	15585 : 1;
	15586 : 1;
	15587 : 1;
	15588 : 1;
	15589 : 1;
	15590 : 1;
	15591 : 1;
	15592 : 1;
	15593 : 1;
	15594 : 1;
	15595 : 1;
	15596 : 1;
	15597 : 1;
	15598 : 1;
	15599 : 1;
	15600 : 1;
	15601 : 1;
	15602 : 1;
	15603 : 1;
	15604 : 1;
	15605 : 1;
	15606 : 1;
	15607 : 1;
	15608 : 1;
	15609 : 1;
	15610 : 1;
	15611 : 1;
	15612 : 1;
	15613 : 1;
	15614 : 1;
	15615 : 1;
	15616 : 1;
	15617 : 1;
	15618 : 1;
	15619 : 1;
	15620 : 1;
	15621 : 1;
	15622 : 1;
	15623 : 1;
	15624 : 1;
	15625 : 1;
	15626 : 1;
	15627 : 1;
	15628 : 1;
	15629 : 1;
	15630 : 1;
	15631 : 1;
	15632 : 1;
	15633 : 1;
	15634 : 1;
	15635 : 1;
	15636 : 1;
	15637 : 1;
	15638 : 1;
	15639 : 1;
	15640 : 1;
	15641 : 1;
	15642 : 1;
	15643 : 1;
	15644 : 1;
	15645 : 1;
	15646 : 1;
	15647 : 1;
	15648 : 1;
	15649 : 1;
	15650 : 1;
	15651 : 1;
	15652 : 1;
	15653 : 1;
	15654 : 1;
	15655 : 1;
	15656 : 1;
	15657 : 1;
	15658 : 1;
	15659 : 1;
	15660 : 1;
	15661 : 1;
	15662 : 1;
	15663 : 1;
	15664 : 1;
	15665 : 1;
	15666 : 1;
	15667 : 1;
	15668 : 1;
	15669 : 1;
	15670 : 1;
	15671 : 1;
	15672 : 1;
	15673 : 1;
	15674 : 1;
	15675 : 1;
	15676 : 1;
	15677 : 1;
	15678 : 1;
	15679 : 1;
	15680 : 1;
	15681 : 1;
	15682 : 1;
	15683 : 1;
	15684 : 1;
	15685 : 1;
	15686 : 1;
	15687 : 1;
	15688 : 1;
	15689 : 1;
	15690 : 1;
	15691 : 1;
	15692 : 1;
	15693 : 1;
	15694 : 1;
	15695 : 1;
	15696 : 1;
	15697 : 1;
	15698 : 1;
	15699 : 1;
	15700 : 1;
	15701 : 1;
	15702 : 1;
	15703 : 1;
	15704 : 1;
	15705 : 1;
	15706 : 1;
	15707 : 1;
	15708 : 1;
	15709 : 1;
	15710 : 1;
	15711 : 1;
	15712 : 1;
	15713 : 1;
	15714 : 1;
	15715 : 1;
	15716 : 1;
	15717 : 1;
	15718 : 1;
	15719 : 1;
	15720 : 1;
	15721 : 1;
	15722 : 1;
	15723 : 1;
	15724 : 1;
	15725 : 1;
	15726 : 1;
	15727 : 1;
	15728 : 1;
	15729 : 1;
	15730 : 1;
	15731 : 1;
	15732 : 1;
	15733 : 1;
	15734 : 1;
	15735 : 1;
	15736 : 1;
	15737 : 1;
	15738 : 1;
	15739 : 1;
	15740 : 1;
	15741 : 1;
	15742 : 1;
	15743 : 1;
	15744 : 1;
	15745 : 1;
	15746 : 1;
	15747 : 1;
	15748 : 1;
	15749 : 1;
	15750 : 1;
	15751 : 1;
	15752 : 1;
	15753 : 1;
	15754 : 1;
	15755 : 1;
	15756 : 1;
	15757 : 1;
	15758 : 1;
	15759 : 1;
	15760 : 1;
	15761 : 1;
	15762 : 1;
	15763 : 1;
	15764 : 1;
	15765 : 1;
	15766 : 1;
	15767 : 1;
	15768 : 1;
	15769 : 1;
	15770 : 1;
	15771 : 1;
	15772 : 1;
	15773 : 1;
	15774 : 1;
	15775 : 1;
	15776 : 1;
	15777 : 1;
	15778 : 1;
	15779 : 1;
	15780 : 1;
	15781 : 1;
	15782 : 1;
	15783 : 1;
	15784 : 1;
	15785 : 1;
	15786 : 1;
	15787 : 1;
	15788 : 1;
	15789 : 1;
	15790 : 1;
	15791 : 1;
	15792 : 1;
	15793 : 1;
	15794 : 1;
	15795 : 1;
	15796 : 1;
	15797 : 1;
	15798 : 1;
	15799 : 1;
	15800 : 1;
	15801 : 1;
	15802 : 1;
	15803 : 1;
	15804 : 1;
	15805 : 1;
	15806 : 1;
	15807 : 1;
	15808 : 1;
	15809 : 1;
	15810 : 1;
	15811 : 1;
	15812 : 1;
	15813 : 1;
	15814 : 1;
	15815 : 1;
	15816 : 1;
	15817 : 1;
	15818 : 1;
	15819 : 1;
	15820 : 1;
	15821 : 1;
	15822 : 1;
	15823 : 1;
	15824 : 1;
	15825 : 1;
	15826 : 1;
	15827 : 1;
	15828 : 1;
	15829 : 1;
	15830 : 1;
	15831 : 1;
	15832 : 1;
	15833 : 1;
	15834 : 1;
	15835 : 1;
	15836 : 1;
	15837 : 1;
	15838 : 1;
	15839 : 1;
	15840 : 1;
	15841 : 1;
	15842 : 1;
	15843 : 1;
	15844 : 1;
	15845 : 1;
	15846 : 1;
	15847 : 1;
	15848 : 1;
	15849 : 1;
	15850 : 1;
	15851 : 1;
	15852 : 1;
	15853 : 1;
	15854 : 1;
	15855 : 1;
	15856 : 1;
	15857 : 1;
	15858 : 1;
	15859 : 1;
	15860 : 1;
	15861 : 1;
	15862 : 1;
	15863 : 1;
	15864 : 1;
	15865 : 1;
	15866 : 1;
	15867 : 1;
	15868 : 1;
	15869 : 1;
	15870 : 1;
	15871 : 1;
	15872 : 1;
	15873 : 1;
	15874 : 1;
	15875 : 1;
	15876 : 1;
	15877 : 1;
	15878 : 1;
	15879 : 1;
	15880 : 1;
	15881 : 1;
	15882 : 1;
	15883 : 1;
	15884 : 1;
	15885 : 1;
	15886 : 1;
	15887 : 1;
	15888 : 1;
	15889 : 1;
	15890 : 1;
	15891 : 1;
	15892 : 1;
	15893 : 1;
	15894 : 1;
	15895 : 1;
	15896 : 1;
	15897 : 1;
	15898 : 1;
	15899 : 1;
	15900 : 1;
	15901 : 1;
	15902 : 1;
	15903 : 1;
	15904 : 1;
	15905 : 1;
	15906 : 1;
	15907 : 1;
	15908 : 1;
	15909 : 1;
	15910 : 1;
	15911 : 1;
	15912 : 1;
	15913 : 1;
	15914 : 1;
	15915 : 1;
	15916 : 1;
	15917 : 1;
	15918 : 1;
	15919 : 1;
	15920 : 1;
	15921 : 1;
	15922 : 1;
	15923 : 1;
	15924 : 1;
	15925 : 1;
	15926 : 1;
	15927 : 1;
	15928 : 1;
	15929 : 1;
	15930 : 1;
	15931 : 1;
	15932 : 1;
	15933 : 1;
	15934 : 1;
	15935 : 1;
	15936 : 1;
	15937 : 1;
	15938 : 1;
	15939 : 1;
	15940 : 1;
	15941 : 1;
	15942 : 1;
	15943 : 1;
	15944 : 1;
	15945 : 1;
	15946 : 1;
	15947 : 1;
	15948 : 1;
	15949 : 1;
	15950 : 1;
	15951 : 1;
	15952 : 1;
	15953 : 1;
	15954 : 1;
	15955 : 1;
	15956 : 1;
	15957 : 1;
	15958 : 1;
	15959 : 1;
	15960 : 1;
	15961 : 1;
	15962 : 1;
	15963 : 1;
	15964 : 1;
	15965 : 1;
	15966 : 1;
	15967 : 1;
	15968 : 1;
	15969 : 1;
	15970 : 1;
	15971 : 1;
	15972 : 1;
	15973 : 1;
	15974 : 1;
	15975 : 1;
	15976 : 1;
	15977 : 1;
	15978 : 1;
	15979 : 1;
	15980 : 1;
	15981 : 1;
	15982 : 1;
	15983 : 1;
	15984 : 1;
	15985 : 1;
	15986 : 1;
	15987 : 1;
	15988 : 1;
	15989 : 1;
	15990 : 1;
	15991 : 1;
	15992 : 1;
	15993 : 1;
	15994 : 1;
	15995 : 1;
	15996 : 1;
	15997 : 1;
	15998 : 1;
	15999 : 1;
	16000 : 1;
	16001 : 1;
	16002 : 1;
	16003 : 1;
	16004 : 1;
	16005 : 1;
	16006 : 1;
	16007 : 1;
	16008 : 1;
	16009 : 1;
	16010 : 1;
	16011 : 1;
	16012 : 1;
	16013 : 1;
	16014 : 1;
	16015 : 1;
	16016 : 1;
	16017 : 1;
	16018 : 1;
	16019 : 1;
	16020 : 1;
	16021 : 1;
	16022 : 1;
	16023 : 1;
	16024 : 1;
	16025 : 1;
	16026 : 1;
	16027 : 1;
	16028 : 1;
	16029 : 1;
	16030 : 1;
	16031 : 1;
	16032 : 1;
	16033 : 1;
	16034 : 1;
	16035 : 1;
	16036 : 1;
	16037 : 1;
	16038 : 1;
	16039 : 1;
	16040 : 1;
	16041 : 1;
	16042 : 1;
	16043 : 1;
	16044 : 1;
	16045 : 1;
	16046 : 1;
	16047 : 1;
	16048 : 1;
	16049 : 1;
	16050 : 1;
	16051 : 1;
	16052 : 1;
	16053 : 1;
	16054 : 1;
	16055 : 1;
	16056 : 1;
	16057 : 1;
	16058 : 1;
	16059 : 1;
	16060 : 1;
	16061 : 1;
	16062 : 1;
	16063 : 1;
	16064 : 1;
	16065 : 1;
	16066 : 1;
	16067 : 1;
	16068 : 1;
	16069 : 1;
	16070 : 1;
	16071 : 1;
	16072 : 1;
	16073 : 1;
	16074 : 1;
	16075 : 1;
	16076 : 1;
	16077 : 1;
	16078 : 1;
	16079 : 1;
	16080 : 1;
	16081 : 1;
	16082 : 1;
	16083 : 1;
	16084 : 1;
	16085 : 1;
	16086 : 1;
	16087 : 1;
	16088 : 1;
	16089 : 1;
	16090 : 1;
	16091 : 1;
	16092 : 1;
	16093 : 1;
	16094 : 1;
	16095 : 1;
	16096 : 1;
	16097 : 1;
	16098 : 1;
	16099 : 1;
	16100 : 1;
	16101 : 1;
	16102 : 1;
	16103 : 1;
	16104 : 1;
	16105 : 1;
	16106 : 1;
	16107 : 1;
	16108 : 1;
	16109 : 1;
	16110 : 1;
	16111 : 1;
	16112 : 1;
	16113 : 1;
	16114 : 1;
	16115 : 1;
	16116 : 1;
	16117 : 1;
	16118 : 1;
	16119 : 1;
	16120 : 1;
	16121 : 1;
	16122 : 1;
	16123 : 1;
	16124 : 1;
	16125 : 1;
	16126 : 1;
	16127 : 1;
	16128 : 1;
	16129 : 1;
	16130 : 1;
	16131 : 1;
	16132 : 1;
	16133 : 1;
	16134 : 1;
	16135 : 1;
	16136 : 1;
	16137 : 1;
	16138 : 1;
	16139 : 1;
	16140 : 1;
	16141 : 1;
	16142 : 1;
	16143 : 1;
	16144 : 1;
	16145 : 1;
	16146 : 1;
	16147 : 1;
	16148 : 1;
	16149 : 1;
	16150 : 1;
	16151 : 1;
	16152 : 1;
	16153 : 1;
	16154 : 1;
	16155 : 1;
	16156 : 1;
	16157 : 1;
	16158 : 1;
	16159 : 1;
	16160 : 1;
	16161 : 1;
	16162 : 1;
	16163 : 1;
	16164 : 1;
	16165 : 1;
	16166 : 1;
	16167 : 1;
	16168 : 1;
	16169 : 1;
	16170 : 1;
	16171 : 1;
	16172 : 1;
	16173 : 1;
	16174 : 1;
	16175 : 1;
	16176 : 1;
	16177 : 1;
	16178 : 1;
	16179 : 1;
	16180 : 1;
	16181 : 1;
	16182 : 1;
	16183 : 1;
	16184 : 1;
	16185 : 1;
	16186 : 1;
	16187 : 1;
	16188 : 1;
	16189 : 1;
	16190 : 1;
	16191 : 1;
	16192 : 1;
	16193 : 1;
	16194 : 1;
	16195 : 1;
	16196 : 1;
	16197 : 1;
	16198 : 1;
	16199 : 1;
	16200 : 1;
	16201 : 1;
	16202 : 1;
	16203 : 1;
	16204 : 1;
	16205 : 1;
	16206 : 1;
	16207 : 1;
	16208 : 1;
	16209 : 1;
	16210 : 1;
	16211 : 1;
	16212 : 1;
	16213 : 1;
	16214 : 1;
	16215 : 1;
	16216 : 1;
	16217 : 1;
	16218 : 1;
	16219 : 1;
	16220 : 1;
	16221 : 1;
	16222 : 1;
	16223 : 1;
	16224 : 1;
	16225 : 1;
	16226 : 1;
	16227 : 1;
	16228 : 1;
	16229 : 1;
	16230 : 1;
	16231 : 1;
	16232 : 1;
	16233 : 1;
	16234 : 1;
	16235 : 1;
	16236 : 1;
	16237 : 1;
	16238 : 1;
	16239 : 1;
	16240 : 1;
	16241 : 1;
	16242 : 1;
	16243 : 1;
	16244 : 1;
	16245 : 1;
	16246 : 1;
	16247 : 1;
	16248 : 1;
	16249 : 1;
	16250 : 1;
	16251 : 1;
	16252 : 1;
	16253 : 1;
	16254 : 1;
	16255 : 1;
	16256 : 1;
	16257 : 1;
	16258 : 1;
	16259 : 1;
	16260 : 1;
	16261 : 1;
	16262 : 1;
	16263 : 1;
	16264 : 1;
	16265 : 1;
	16266 : 1;
	16267 : 1;
	16268 : 1;
	16269 : 1;
	16270 : 1;
	16271 : 1;
	16272 : 1;
	16273 : 1;
	16274 : 1;
	16275 : 1;
	16276 : 1;
	16277 : 1;
	16278 : 1;
	16279 : 1;
	16280 : 1;
	16281 : 1;
	16282 : 1;
	16283 : 1;
	16284 : 1;
	16285 : 1;
	16286 : 1;
	16287 : 1;
	16288 : 1;
	16289 : 1;
	16290 : 1;
	16291 : 1;
	16292 : 1;
	16293 : 1;
	16294 : 1;
	16295 : 1;
	16296 : 1;
	16297 : 1;
	16298 : 1;
	16299 : 1;
	16300 : 1;
	16301 : 1;
	16302 : 1;
	16303 : 1;
	16304 : 1;
	16305 : 1;
	16306 : 1;
	16307 : 1;
	16308 : 1;
	16309 : 1;
	16310 : 1;
	16311 : 1;
	16312 : 1;
	16313 : 1;
	16314 : 1;
	16315 : 1;
	16316 : 1;
	16317 : 1;
	16318 : 1;
	16319 : 1;
	16320 : 1;
	16321 : 1;
	16322 : 1;
	16323 : 1;
	16324 : 1;
	16325 : 1;
	16326 : 1;
	16327 : 1;
	16328 : 1;
	16329 : 1;
	16330 : 1;
	16331 : 1;
	16332 : 1;
	16333 : 1;
	16334 : 1;
	16335 : 1;
	16336 : 1;
	16337 : 1;
	16338 : 1;
	16339 : 1;
	16340 : 1;
	16341 : 1;
	16342 : 1;
	16343 : 1;
	16344 : 1;
	16345 : 1;
	16346 : 1;
	16347 : 1;
	16348 : 1;
	16349 : 1;
	16350 : 1;
	16351 : 1;
	16352 : 1;
	16353 : 1;
	16354 : 1;
	16355 : 1;
	16356 : 1;
	16357 : 1;
	16358 : 1;
	16359 : 1;
	16360 : 1;
	16361 : 1;
	16362 : 1;
	16363 : 1;
	16364 : 1;
	16365 : 1;
	16366 : 1;
	16367 : 1;
	16368 : 1;
	16369 : 1;
	16370 : 1;
	16371 : 1;
	16372 : 1;
	16373 : 1;
	16374 : 1;
	16375 : 1;
	16376 : 1;
	16377 : 1;
	16378 : 1;
	16379 : 1;
	16380 : 1;
	16381 : 1;
	16382 : 1;
	16383 : 1;
	16384 : 1;
	16385 : 1;
	16386 : 1;
	16387 : 1;
	16388 : 1;
	16389 : 1;
	16390 : 1;
	16391 : 1;
	16392 : 1;
	16393 : 1;
	16394 : 1;
	16395 : 1;
	16396 : 1;
	16397 : 1;
	16398 : 1;
	16399 : 1;
	16400 : 1;
	16401 : 1;
	16402 : 1;
	16403 : 1;
	16404 : 1;
	16405 : 1;
	16406 : 1;
	16407 : 1;
	16408 : 1;
	16409 : 1;
	16410 : 1;
	16411 : 1;
	16412 : 1;
	16413 : 1;
	16414 : 1;
	16415 : 1;
	16416 : 1;
	16417 : 1;
	16418 : 1;
	16419 : 1;
	16420 : 1;
	16421 : 1;
	16422 : 1;
	16423 : 1;
	16424 : 1;
	16425 : 1;
	16426 : 1;
	16427 : 1;
	16428 : 1;
	16429 : 1;
	16430 : 1;
	16431 : 1;
	16432 : 1;
	16433 : 1;
	16434 : 1;
	16435 : 1;
	16436 : 1;
	16437 : 1;
	16438 : 1;
	16439 : 1;
	16440 : 1;
	16441 : 1;
	16442 : 1;
	16443 : 1;
	16444 : 1;
	16445 : 1;
	16446 : 1;
	16447 : 1;
	16448 : 1;
	16449 : 1;
	16450 : 1;
	16451 : 1;
	16452 : 1;
	16453 : 1;
	16454 : 1;
	16455 : 1;
	16456 : 1;
	16457 : 1;
	16458 : 1;
	16459 : 1;
	16460 : 1;
	16461 : 1;
	16462 : 1;
	16463 : 1;
	16464 : 1;
	16465 : 1;
	16466 : 1;
	16467 : 1;
	16468 : 1;
	16469 : 1;
	16470 : 1;
	16471 : 1;
	16472 : 1;
	16473 : 1;
	16474 : 1;
	16475 : 1;
	16476 : 1;
	16477 : 1;
	16478 : 1;
	16479 : 1;
	16480 : 1;
	16481 : 1;
	16482 : 1;
	16483 : 1;
	16484 : 1;
	16485 : 1;
	16486 : 1;
	16487 : 1;
	16488 : 1;
	16489 : 1;
	16490 : 1;
	16491 : 1;
	16492 : 1;
	16493 : 1;
	16494 : 1;
	16495 : 1;
	16496 : 1;
	16497 : 1;
	16498 : 1;
	16499 : 1;
	16500 : 1;
	16501 : 1;
	16502 : 1;
	16503 : 1;
	16504 : 1;
	16505 : 1;
	16506 : 1;
	16507 : 1;
	16508 : 1;
	16509 : 1;
	16510 : 1;
	16511 : 1;
	16512 : 1;
	16513 : 1;
	16514 : 1;
	16515 : 1;
	16516 : 1;
	16517 : 1;
	16518 : 1;
	16519 : 1;
	16520 : 1;
	16521 : 1;
	16522 : 1;
	16523 : 1;
	16524 : 1;
	16525 : 1;
	16526 : 1;
	16527 : 1;
	16528 : 1;
	16529 : 1;
	16530 : 1;
	16531 : 1;
	16532 : 1;
	16533 : 1;
	16534 : 1;
	16535 : 1;
	16536 : 1;
	16537 : 1;
	16538 : 1;
	16539 : 1;
	16540 : 1;
	16541 : 1;
	16542 : 1;
	16543 : 1;
	16544 : 1;
	16545 : 1;
	16546 : 1;
	16547 : 1;
	16548 : 1;
	16549 : 1;
	16550 : 1;
	16551 : 1;
	16552 : 1;
	16553 : 1;
	16554 : 1;
	16555 : 1;
	16556 : 1;
	16557 : 1;
	16558 : 1;
	16559 : 1;
	16560 : 1;
	16561 : 1;
	16562 : 1;
	16563 : 1;
	16564 : 1;
	16565 : 1;
	16566 : 1;
	16567 : 1;
	16568 : 1;
	16569 : 1;
	16570 : 1;
	16571 : 1;
	16572 : 1;
	16573 : 1;
	16574 : 1;
	16575 : 1;
	16576 : 1;
	16577 : 1;
	16578 : 1;
	16579 : 1;
	16580 : 1;
	16581 : 1;
	16582 : 1;
	16583 : 1;
	16584 : 1;
	16585 : 1;
	16586 : 1;
	16587 : 1;
	16588 : 1;
	16589 : 1;
	16590 : 1;
	16591 : 1;
	16592 : 1;
	16593 : 1;
	16594 : 1;
	16595 : 1;
	16596 : 1;
	16597 : 1;
	16598 : 1;
	16599 : 1;
	16600 : 1;
	16601 : 1;
	16602 : 1;
	16603 : 1;
	16604 : 1;
	16605 : 1;
	16606 : 1;
	16607 : 1;
	16608 : 1;
	16609 : 1;
	16610 : 1;
	16611 : 1;
	16612 : 1;
	16613 : 1;
	16614 : 1;
	16615 : 1;
	16616 : 1;
	16617 : 1;
	16618 : 1;
	16619 : 1;
	16620 : 1;
	16621 : 1;
	16622 : 1;
	16623 : 1;
	16624 : 1;
	16625 : 1;
	16626 : 1;
	16627 : 1;
	16628 : 1;
	16629 : 1;
	16630 : 1;
	16631 : 1;
	16632 : 1;
	16633 : 1;
	16634 : 1;
	16635 : 1;
	16636 : 1;
	16637 : 1;
	16638 : 1;
	16639 : 1;
	16640 : 1;
	16641 : 1;
	16642 : 1;
	16643 : 1;
	16644 : 1;
	16645 : 1;
	16646 : 1;
	16647 : 1;
	16648 : 1;
	16649 : 1;
	16650 : 1;
	16651 : 1;
	16652 : 1;
	16653 : 1;
	16654 : 1;
	16655 : 1;
	16656 : 1;
	16657 : 1;
	16658 : 1;
	16659 : 1;
	16660 : 1;
	16661 : 1;
	16662 : 1;
	16663 : 1;
	16664 : 1;
	16665 : 1;
	16666 : 1;
	16667 : 1;
	16668 : 1;
	16669 : 1;
	16670 : 1;
	16671 : 1;
	16672 : 1;
	16673 : 1;
	16674 : 1;
	16675 : 1;
	16676 : 1;
	16677 : 1;
	16678 : 1;
	16679 : 1;
	16680 : 1;
	16681 : 1;
	16682 : 1;
	16683 : 1;
	16684 : 1;
	16685 : 1;
	16686 : 1;
	16687 : 1;
	16688 : 1;
	16689 : 1;
	16690 : 1;
	16691 : 1;
	16692 : 1;
	16693 : 1;
	16694 : 1;
	16695 : 1;
	16696 : 1;
	16697 : 1;
	16698 : 1;
	16699 : 1;
	16700 : 1;
	16701 : 1;
	16702 : 1;
	16703 : 1;
	16704 : 1;
	16705 : 1;
	16706 : 1;
	16707 : 1;
	16708 : 1;
	16709 : 1;
	16710 : 1;
	16711 : 1;
	16712 : 1;
	16713 : 1;
	16714 : 1;
	16715 : 1;
	16716 : 1;
	16717 : 1;
	16718 : 1;
	16719 : 1;
	16720 : 1;
	16721 : 1;
	16722 : 1;
	16723 : 1;
	16724 : 1;
	16725 : 1;
	16726 : 1;
	16727 : 1;
	16728 : 1;
	16729 : 1;
	16730 : 1;
	16731 : 1;
	16732 : 1;
	16733 : 1;
	16734 : 1;
	16735 : 1;
	16736 : 1;
	16737 : 1;
	16738 : 1;
	16739 : 1;
	16740 : 1;
	16741 : 1;
	16742 : 1;
	16743 : 1;
	16744 : 1;
	16745 : 1;
	16746 : 1;
	16747 : 1;
	16748 : 1;
	16749 : 1;
	16750 : 1;
	16751 : 1;
	16752 : 1;
	16753 : 1;
	16754 : 1;
	16755 : 1;
	16756 : 1;
	16757 : 1;
	16758 : 1;
	16759 : 1;
	16760 : 1;
	16761 : 1;
	16762 : 1;
	16763 : 1;
	16764 : 1;
	16765 : 1;
	16766 : 1;
	16767 : 1;
	16768 : 1;
	16769 : 1;
	16770 : 1;
	16771 : 1;
	16772 : 1;
	16773 : 1;
	16774 : 1;
	16775 : 1;
	16776 : 1;
	16777 : 1;
	16778 : 1;
	16779 : 1;
	16780 : 1;
	16781 : 1;
	16782 : 1;
	16783 : 1;
	16784 : 1;
	16785 : 1;
	16786 : 1;
	16787 : 1;
	16788 : 1;
	16789 : 1;
	16790 : 1;
	16791 : 1;
	16792 : 1;
	16793 : 1;
	16794 : 1;
	16795 : 1;
	16796 : 1;
	16797 : 1;
	16798 : 1;
	16799 : 1;
	16800 : 1;
	16801 : 1;
	16802 : 1;
	16803 : 1;
	16804 : 1;
	16805 : 1;
	16806 : 1;
	16807 : 1;
	16808 : 1;
	16809 : 1;
	16810 : 1;
	16811 : 1;
	16812 : 1;
	16813 : 1;
	16814 : 1;
	16815 : 1;
	16816 : 1;
	16817 : 1;
	16818 : 1;
	16819 : 1;
	16820 : 1;
	16821 : 1;
	16822 : 1;
	16823 : 1;
	16824 : 1;
	16825 : 1;
	16826 : 1;
	16827 : 1;
	16828 : 1;
	16829 : 1;
	16830 : 1;
	16831 : 1;
	16832 : 1;
	16833 : 1;
	16834 : 1;
	16835 : 1;
	16836 : 1;
	16837 : 1;
	16838 : 1;
	16839 : 1;
	16840 : 1;
	16841 : 1;
	16842 : 1;
	16843 : 1;
	16844 : 1;
	16845 : 1;
	16846 : 1;
	16847 : 1;
	16848 : 1;
	16849 : 1;
	16850 : 1;
	16851 : 1;
	16852 : 1;
	16853 : 1;
	16854 : 1;
	16855 : 1;
	16856 : 1;
	16857 : 1;
	16858 : 1;
	16859 : 1;
	16860 : 1;
	16861 : 1;
	16862 : 1;
	16863 : 1;
	16864 : 1;
	16865 : 1;
	16866 : 1;
	16867 : 1;
	16868 : 1;
	16869 : 1;
	16870 : 1;
	16871 : 1;
	16872 : 1;
	16873 : 1;
	16874 : 1;
	16875 : 1;
	16876 : 1;
	16877 : 1;
	16878 : 1;
	16879 : 1;
	16880 : 1;
	16881 : 1;
	16882 : 1;
	16883 : 1;
	16884 : 1;
	16885 : 1;
	16886 : 1;
	16887 : 1;
	16888 : 1;
	16889 : 1;
	16890 : 1;
	16891 : 1;
	16892 : 1;
	16893 : 1;
	16894 : 1;
	16895 : 1;
	16896 : 1;
	16897 : 1;
	16898 : 1;
	16899 : 1;
	16900 : 1;
	16901 : 1;
	16902 : 1;
	16903 : 1;
	16904 : 1;
	16905 : 1;
	16906 : 1;
	16907 : 1;
	16908 : 1;
	16909 : 1;
	16910 : 1;
	16911 : 1;
	16912 : 1;
	16913 : 1;
	16914 : 1;
	16915 : 1;
	16916 : 1;
	16917 : 1;
	16918 : 1;
	16919 : 1;
	16920 : 1;
	16921 : 1;
	16922 : 1;
	16923 : 1;
	16924 : 1;
	16925 : 1;
	16926 : 1;
	16927 : 1;
	16928 : 1;
	16929 : 1;
	16930 : 1;
	16931 : 1;
	16932 : 1;
	16933 : 1;
	16934 : 1;
	16935 : 1;
	16936 : 1;
	16937 : 1;
	16938 : 1;
	16939 : 1;
	16940 : 1;
	16941 : 1;
	16942 : 1;
	16943 : 1;
	16944 : 1;
	16945 : 1;
	16946 : 1;
	16947 : 1;
	16948 : 1;
	16949 : 1;
	16950 : 1;
	16951 : 1;
	16952 : 1;
	16953 : 1;
	16954 : 1;
	16955 : 1;
	16956 : 1;
	16957 : 1;
	16958 : 1;
	16959 : 1;
	16960 : 1;
	16961 : 1;
	16962 : 1;
	16963 : 1;
	16964 : 1;
	16965 : 1;
	16966 : 1;
	16967 : 1;
	16968 : 1;
	16969 : 1;
	16970 : 1;
	16971 : 1;
	16972 : 1;
	16973 : 1;
	16974 : 1;
	16975 : 1;
	16976 : 1;
	16977 : 1;
	16978 : 1;
	16979 : 1;
	16980 : 1;
	16981 : 1;
	16982 : 1;
	16983 : 1;
	16984 : 1;
	16985 : 1;
	16986 : 1;
	16987 : 1;
	16988 : 1;
	16989 : 1;
	16990 : 1;
	16991 : 1;
	16992 : 1;
	16993 : 1;
	16994 : 1;
	16995 : 1;
	16996 : 1;
	16997 : 1;
	16998 : 1;
	16999 : 1;
	17000 : 1;
	17001 : 1;
	17002 : 1;
	17003 : 1;
	17004 : 1;
	17005 : 1;
	17006 : 1;
	17007 : 1;
	17008 : 1;
	17009 : 1;
	17010 : 1;
	17011 : 1;
	17012 : 1;
	17013 : 1;
	17014 : 1;
	17015 : 1;
	17016 : 1;
	17017 : 1;
	17018 : 1;
	17019 : 1;
	17020 : 1;
	17021 : 1;
	17022 : 1;
	17023 : 1;
	17024 : 1;
	17025 : 1;
	17026 : 1;
	17027 : 1;
	17028 : 1;
	17029 : 1;
	17030 : 1;
	17031 : 1;
	17032 : 1;
	17033 : 1;
	17034 : 1;
	17035 : 1;
	17036 : 1;
	17037 : 1;
	17038 : 1;
	17039 : 1;
	17040 : 1;
	17041 : 1;
	17042 : 1;
	17043 : 1;
	17044 : 1;
	17045 : 1;
	17046 : 1;
	17047 : 1;
	17048 : 1;
	17049 : 1;
	17050 : 0;
	17051 : 0;
	17052 : 0;
	17053 : 0;
	17054 : 1;
	17055 : 1;
	17056 : 0;
	17057 : 0;
	17058 : 0;
	17059 : 0;
	17060 : 1;
	17061 : 1;
	17062 : 1;
	17063 : 1;
	17064 : 0;
	17065 : 0;
	17066 : 0;
	17067 : 0;
	17068 : 1;
	17069 : 1;
	17070 : 1;
	17071 : 1;
	17072 : 1;
	17073 : 1;
	17074 : 1;
	17075 : 1;
	17076 : 1;
	17077 : 1;
	17078 : 1;
	17079 : 1;
	17080 : 1;
	17081 : 1;
	17082 : 1;
	17083 : 1;
	17084 : 1;
	17085 : 1;
	17086 : 0;
	17087 : 0;
	17088 : 1;
	17089 : 1;
	17090 : 1;
	17091 : 1;
	17092 : 1;
	17093 : 1;
	17094 : 1;
	17095 : 1;
	17096 : 1;
	17097 : 1;
	17098 : 1;
	17099 : 1;
	17100 : 1;
	17101 : 1;
	17102 : 1;
	17103 : 1;
	17104 : 1;
	17105 : 1;
	17106 : 1;
	17107 : 1;
	17108 : 1;
	17109 : 1;
	17110 : 1;
	17111 : 0;
	17112 : 0;
	17113 : 0;
	17114 : 0;
	17115 : 1;
	17116 : 1;
	17117 : 0;
	17118 : 0;
	17119 : 0;
	17120 : 0;
	17121 : 1;
	17122 : 1;
	17123 : 1;
	17124 : 1;
	17125 : 0;
	17126 : 0;
	17127 : 0;
	17128 : 0;
	17129 : 0;
	17130 : 1;
	17131 : 1;
	17132 : 1;
	17133 : 1;
	17134 : 1;
	17135 : 1;
	17136 : 1;
	17137 : 1;
	17138 : 1;
	17139 : 1;
	17140 : 1;
	17141 : 1;
	17142 : 1;
	17143 : 1;
	17144 : 1;
	17145 : 1;
	17146 : 1;
	17147 : 1;
	17148 : 1;
	17149 : 1;
	17150 : 1;
	17151 : 1;
	17152 : 1;
	17153 : 1;
	17154 : 1;
	17155 : 1;
	17156 : 1;
	17157 : 1;
	17158 : 1;
	17159 : 1;
	17160 : 1;
	17161 : 1;
	17162 : 1;
	17163 : 0;
	17164 : 0;
	17165 : 1;
	17166 : 1;
	17167 : 1;
	17168 : 1;
	17169 : 1;
	17170 : 1;
	17171 : 1;
	17172 : 1;
	17173 : 1;
	17174 : 1;
	17175 : 1;
	17176 : 1;
	17177 : 1;
	17178 : 1;
	17179 : 1;
	17180 : 1;
	17181 : 1;
	17182 : 1;
	17183 : 1;
	17184 : 1;
	17185 : 1;
	17186 : 1;
	17187 : 1;
	17188 : 1;
	17189 : 1;
	17190 : 1;
	17191 : 1;
	17192 : 1;
	17193 : 1;
	17194 : 1;
	17195 : 1;
	17196 : 1;
	17197 : 1;
	17198 : 1;
	17199 : 1;
	17200 : 1;
	17201 : 1;
	17202 : 1;
	17203 : 1;
	17204 : 1;
	17205 : 1;
	17206 : 1;
	17207 : 1;
	17208 : 1;
	17209 : 1;
	17210 : 1;
	17211 : 1;
	17212 : 1;
	17213 : 1;
	17214 : 1;
	17215 : 1;
	17216 : 1;
	17217 : 1;
	17218 : 1;
	17219 : 1;
	17220 : 1;
	17221 : 1;
	17222 : 1;
	17223 : 1;
	17224 : 0;
	17225 : 1;
	17226 : 1;
	17227 : 1;
	17228 : 1;
	17229 : 1;
	17230 : 1;
	17231 : 1;
	17232 : 1;
	17233 : 1;
	17234 : 1;
	17235 : 1;
	17236 : 1;
	17237 : 1;
	17238 : 0;
	17239 : 0;
	17240 : 1;
	17241 : 1;
	17242 : 1;
	17243 : 1;
	17244 : 1;
	17245 : 1;
	17246 : 1;
	17247 : 1;
	17248 : 1;
	17249 : 1;
	17250 : 1;
	17251 : 0;
	17252 : 0;
	17253 : 1;
	17254 : 1;
	17255 : 1;
	17256 : 1;
	17257 : 1;
	17258 : 1;
	17259 : 1;
	17260 : 1;
	17261 : 1;
	17262 : 1;
	17263 : 1;
	17264 : 1;
	17265 : 1;
	17266 : 1;
	17267 : 1;
	17268 : 1;
	17269 : 1;
	17270 : 1;
	17271 : 0;
	17272 : 1;
	17273 : 1;
	17274 : 1;
	17275 : 1;
	17276 : 1;
	17277 : 1;
	17278 : 1;
	17279 : 1;
	17280 : 1;
	17281 : 1;
	17282 : 1;
	17283 : 1;
	17284 : 1;
	17285 : 1;
	17286 : 1;
	17287 : 1;
	17288 : 1;
	17289 : 0;
	17290 : 1;
	17291 : 1;
	17292 : 1;
	17293 : 0;
	17294 : 1;
	17295 : 0;
	17296 : 1;
	17297 : 1;
	17298 : 1;
	17299 : 0;
	17300 : 0;
	17301 : 1;
	17302 : 1;
	17303 : 0;
	17304 : 0;
	17305 : 1;
	17306 : 1;
	17307 : 1;
	17308 : 0;
	17309 : 1;
	17310 : 1;
	17311 : 1;
	17312 : 1;
	17313 : 1;
	17314 : 1;
	17315 : 1;
	17316 : 1;
	17317 : 1;
	17318 : 1;
	17319 : 1;
	17320 : 1;
	17321 : 1;
	17322 : 1;
	17323 : 1;
	17324 : 1;
	17325 : 1;
	17326 : 0;
	17327 : 0;
	17328 : 1;
	17329 : 1;
	17330 : 1;
	17331 : 1;
	17332 : 1;
	17333 : 1;
	17334 : 1;
	17335 : 1;
	17336 : 1;
	17337 : 1;
	17338 : 1;
	17339 : 1;
	17340 : 1;
	17341 : 1;
	17342 : 1;
	17343 : 1;
	17344 : 1;
	17345 : 1;
	17346 : 1;
	17347 : 1;
	17348 : 1;
	17349 : 1;
	17350 : 0;
	17351 : 1;
	17352 : 1;
	17353 : 1;
	17354 : 1;
	17355 : 1;
	17356 : 0;
	17357 : 0;
	17358 : 1;
	17359 : 1;
	17360 : 1;
	17361 : 0;
	17362 : 1;
	17363 : 1;
	17364 : 1;
	17365 : 1;
	17366 : 1;
	17367 : 0;
	17368 : 1;
	17369 : 1;
	17370 : 1;
	17371 : 1;
	17372 : 1;
	17373 : 1;
	17374 : 1;
	17375 : 1;
	17376 : 1;
	17377 : 1;
	17378 : 1;
	17379 : 1;
	17380 : 1;
	17381 : 1;
	17382 : 1;
	17383 : 1;
	17384 : 1;
	17385 : 1;
	17386 : 1;
	17387 : 1;
	17388 : 1;
	17389 : 1;
	17390 : 1;
	17391 : 1;
	17392 : 1;
	17393 : 1;
	17394 : 1;
	17395 : 1;
	17396 : 1;
	17397 : 1;
	17398 : 1;
	17399 : 1;
	17400 : 1;
	17401 : 1;
	17402 : 1;
	17403 : 0;
	17404 : 0;
	17405 : 1;
	17406 : 1;
	17407 : 1;
	17408 : 1;
	17409 : 1;
	17410 : 1;
	17411 : 1;
	17412 : 1;
	17413 : 1;
	17414 : 1;
	17415 : 1;
	17416 : 1;
	17417 : 1;
	17418 : 1;
	17419 : 1;
	17420 : 1;
	17421 : 1;
	17422 : 1;
	17423 : 1;
	17424 : 1;
	17425 : 1;
	17426 : 1;
	17427 : 1;
	17428 : 1;
	17429 : 1;
	17430 : 1;
	17431 : 1;
	17432 : 1;
	17433 : 1;
	17434 : 1;
	17435 : 1;
	17436 : 1;
	17437 : 1;
	17438 : 1;
	17439 : 1;
	17440 : 1;
	17441 : 1;
	17442 : 1;
	17443 : 1;
	17444 : 1;
	17445 : 1;
	17446 : 1;
	17447 : 1;
	17448 : 1;
	17449 : 1;
	17450 : 1;
	17451 : 1;
	17452 : 1;
	17453 : 1;
	17454 : 1;
	17455 : 1;
	17456 : 1;
	17457 : 1;
	17458 : 1;
	17459 : 1;
	17460 : 1;
	17461 : 1;
	17462 : 1;
	17463 : 1;
	17464 : 0;
	17465 : 1;
	17466 : 1;
	17467 : 1;
	17468 : 1;
	17469 : 1;
	17470 : 1;
	17471 : 1;
	17472 : 1;
	17473 : 1;
	17474 : 1;
	17475 : 1;
	17476 : 1;
	17477 : 1;
	17478 : 0;
	17479 : 0;
	17480 : 1;
	17481 : 1;
	17482 : 1;
	17483 : 1;
	17484 : 1;
	17485 : 1;
	17486 : 1;
	17487 : 1;
	17488 : 1;
	17489 : 1;
	17490 : 1;
	17491 : 1;
	17492 : 0;
	17493 : 1;
	17494 : 1;
	17495 : 1;
	17496 : 1;
	17497 : 1;
	17498 : 1;
	17499 : 1;
	17500 : 1;
	17501 : 1;
	17502 : 1;
	17503 : 1;
	17504 : 1;
	17505 : 1;
	17506 : 1;
	17507 : 1;
	17508 : 1;
	17509 : 1;
	17510 : 1;
	17511 : 0;
	17512 : 1;
	17513 : 1;
	17514 : 1;
	17515 : 1;
	17516 : 1;
	17517 : 1;
	17518 : 1;
	17519 : 1;
	17520 : 1;
	17521 : 1;
	17522 : 1;
	17523 : 1;
	17524 : 1;
	17525 : 1;
	17526 : 1;
	17527 : 1;
	17528 : 1;
	17529 : 0;
	17530 : 1;
	17531 : 1;
	17532 : 1;
	17533 : 1;
	17534 : 1;
	17535 : 0;
	17536 : 1;
	17537 : 1;
	17538 : 1;
	17539 : 0;
	17540 : 0;
	17541 : 1;
	17542 : 1;
	17543 : 0;
	17544 : 0;
	17545 : 1;
	17546 : 1;
	17547 : 1;
	17548 : 0;
	17549 : 1;
	17550 : 1;
	17551 : 1;
	17552 : 1;
	17553 : 1;
	17554 : 1;
	17555 : 1;
	17556 : 1;
	17557 : 1;
	17558 : 1;
	17559 : 1;
	17560 : 1;
	17561 : 1;
	17562 : 1;
	17563 : 1;
	17564 : 1;
	17565 : 1;
	17566 : 0;
	17567 : 0;
	17568 : 1;
	17569 : 1;
	17570 : 1;
	17571 : 1;
	17572 : 1;
	17573 : 1;
	17574 : 1;
	17575 : 1;
	17576 : 1;
	17577 : 1;
	17578 : 1;
	17579 : 1;
	17580 : 1;
	17581 : 1;
	17582 : 1;
	17583 : 1;
	17584 : 1;
	17585 : 1;
	17586 : 1;
	17587 : 1;
	17588 : 1;
	17589 : 1;
	17590 : 0;
	17591 : 1;
	17592 : 1;
	17593 : 1;
	17594 : 1;
	17595 : 1;
	17596 : 0;
	17597 : 0;
	17598 : 1;
	17599 : 1;
	17600 : 1;
	17601 : 0;
	17602 : 1;
	17603 : 1;
	17604 : 1;
	17605 : 1;
	17606 : 1;
	17607 : 0;
	17608 : 1;
	17609 : 1;
	17610 : 1;
	17611 : 1;
	17612 : 1;
	17613 : 1;
	17614 : 1;
	17615 : 1;
	17616 : 1;
	17617 : 1;
	17618 : 1;
	17619 : 1;
	17620 : 1;
	17621 : 1;
	17622 : 1;
	17623 : 1;
	17624 : 1;
	17625 : 1;
	17626 : 1;
	17627 : 1;
	17628 : 1;
	17629 : 1;
	17630 : 1;
	17631 : 1;
	17632 : 1;
	17633 : 1;
	17634 : 1;
	17635 : 1;
	17636 : 1;
	17637 : 1;
	17638 : 1;
	17639 : 1;
	17640 : 1;
	17641 : 1;
	17642 : 1;
	17643 : 0;
	17644 : 0;
	17645 : 1;
	17646 : 1;
	17647 : 1;
	17648 : 1;
	17649 : 1;
	17650 : 1;
	17651 : 1;
	17652 : 1;
	17653 : 1;
	17654 : 1;
	17655 : 1;
	17656 : 1;
	17657 : 1;
	17658 : 1;
	17659 : 1;
	17660 : 1;
	17661 : 1;
	17662 : 1;
	17663 : 1;
	17664 : 1;
	17665 : 1;
	17666 : 1;
	17667 : 1;
	17668 : 1;
	17669 : 1;
	17670 : 1;
	17671 : 1;
	17672 : 1;
	17673 : 1;
	17674 : 1;
	17675 : 1;
	17676 : 1;
	17677 : 1;
	17678 : 1;
	17679 : 1;
	17680 : 1;
	17681 : 1;
	17682 : 1;
	17683 : 1;
	17684 : 1;
	17685 : 1;
	17686 : 1;
	17687 : 1;
	17688 : 1;
	17689 : 1;
	17690 : 1;
	17691 : 1;
	17692 : 1;
	17693 : 1;
	17694 : 1;
	17695 : 1;
	17696 : 1;
	17697 : 1;
	17698 : 1;
	17699 : 1;
	17700 : 1;
	17701 : 1;
	17702 : 1;
	17703 : 1;
	17704 : 0;
	17705 : 1;
	17706 : 1;
	17707 : 1;
	17708 : 1;
	17709 : 1;
	17710 : 1;
	17711 : 1;
	17712 : 1;
	17713 : 1;
	17714 : 1;
	17715 : 1;
	17716 : 1;
	17717 : 1;
	17718 : 0;
	17719 : 0;
	17720 : 1;
	17721 : 1;
	17722 : 1;
	17723 : 1;
	17724 : 1;
	17725 : 1;
	17726 : 1;
	17727 : 1;
	17728 : 1;
	17729 : 1;
	17730 : 1;
	17731 : 1;
	17732 : 0;
	17733 : 1;
	17734 : 1;
	17735 : 1;
	17736 : 1;
	17737 : 1;
	17738 : 1;
	17739 : 1;
	17740 : 1;
	17741 : 1;
	17742 : 1;
	17743 : 1;
	17744 : 1;
	17745 : 1;
	17746 : 1;
	17747 : 1;
	17748 : 1;
	17749 : 1;
	17750 : 0;
	17751 : 0;
	17752 : 1;
	17753 : 1;
	17754 : 1;
	17755 : 1;
	17756 : 1;
	17757 : 1;
	17758 : 1;
	17759 : 1;
	17760 : 1;
	17761 : 1;
	17762 : 1;
	17763 : 1;
	17764 : 1;
	17765 : 1;
	17766 : 1;
	17767 : 1;
	17768 : 1;
	17769 : 0;
	17770 : 1;
	17771 : 1;
	17772 : 1;
	17773 : 1;
	17774 : 1;
	17775 : 0;
	17776 : 0;
	17777 : 1;
	17778 : 1;
	17779 : 0;
	17780 : 0;
	17781 : 1;
	17782 : 1;
	17783 : 0;
	17784 : 0;
	17785 : 1;
	17786 : 1;
	17787 : 0;
	17788 : 0;
	17789 : 1;
	17790 : 0;
	17791 : 0;
	17792 : 0;
	17793 : 1;
	17794 : 1;
	17795 : 0;
	17796 : 1;
	17797 : 1;
	17798 : 0;
	17799 : 1;
	17800 : 1;
	17801 : 0;
	17802 : 0;
	17803 : 0;
	17804 : 0;
	17805 : 1;
	17806 : 0;
	17807 : 0;
	17808 : 0;
	17809 : 0;
	17810 : 0;
	17811 : 1;
	17812 : 1;
	17813 : 0;
	17814 : 1;
	17815 : 1;
	17816 : 1;
	17817 : 0;
	17818 : 1;
	17819 : 1;
	17820 : 0;
	17821 : 0;
	17822 : 0;
	17823 : 0;
	17824 : 1;
	17825 : 1;
	17826 : 1;
	17827 : 1;
	17828 : 1;
	17829 : 1;
	17830 : 0;
	17831 : 1;
	17832 : 1;
	17833 : 1;
	17834 : 1;
	17835 : 1;
	17836 : 0;
	17837 : 0;
	17838 : 1;
	17839 : 1;
	17840 : 0;
	17841 : 0;
	17842 : 1;
	17843 : 1;
	17844 : 1;
	17845 : 1;
	17846 : 1;
	17847 : 0;
	17848 : 1;
	17849 : 1;
	17850 : 1;
	17851 : 1;
	17852 : 0;
	17853 : 0;
	17854 : 0;
	17855 : 0;
	17856 : 0;
	17857 : 0;
	17858 : 0;
	17859 : 0;
	17860 : 0;
	17861 : 1;
	17862 : 1;
	17863 : 1;
	17864 : 1;
	17865 : 1;
	17866 : 1;
	17867 : 1;
	17868 : 0;
	17869 : 0;
	17870 : 0;
	17871 : 0;
	17872 : 0;
	17873 : 1;
	17874 : 0;
	17875 : 0;
	17876 : 0;
	17877 : 0;
	17878 : 1;
	17879 : 1;
	17880 : 0;
	17881 : 0;
	17882 : 0;
	17883 : 0;
	17884 : 0;
	17885 : 1;
	17886 : 1;
	17887 : 1;
	17888 : 0;
	17889 : 0;
	17890 : 0;
	17891 : 0;
	17892 : 1;
	17893 : 1;
	17894 : 0;
	17895 : 1;
	17896 : 1;
	17897 : 1;
	17898 : 0;
	17899 : 1;
	17900 : 1;
	17901 : 0;
	17902 : 0;
	17903 : 0;
	17904 : 0;
	17905 : 1;
	17906 : 0;
	17907 : 0;
	17908 : 0;
	17909 : 0;
	17910 : 0;
	17911 : 0;
	17912 : 0;
	17913 : 1;
	17914 : 1;
	17915 : 1;
	17916 : 0;
	17917 : 1;
	17918 : 0;
	17919 : 0;
	17920 : 0;
	17921 : 0;
	17922 : 1;
	17923 : 1;
	17924 : 0;
	17925 : 0;
	17926 : 0;
	17927 : 0;
	17928 : 1;
	17929 : 1;
	17930 : 0;
	17931 : 0;
	17932 : 0;
	17933 : 0;
	17934 : 1;
	17935 : 1;
	17936 : 1;
	17937 : 1;
	17938 : 0;
	17939 : 1;
	17940 : 0;
	17941 : 1;
	17942 : 0;
	17943 : 1;
	17944 : 0;
	17945 : 0;
	17946 : 0;
	17947 : 0;
	17948 : 0;
	17949 : 1;
	17950 : 1;
	17951 : 0;
	17952 : 0;
	17953 : 0;
	17954 : 0;
	17955 : 1;
	17956 : 1;
	17957 : 1;
	17958 : 0;
	17959 : 0;
	17960 : 0;
	17961 : 0;
	17962 : 0;
	17963 : 1;
	17964 : 1;
	17965 : 0;
	17966 : 0;
	17967 : 0;
	17968 : 0;
	17969 : 1;
	17970 : 1;
	17971 : 1;
	17972 : 0;
	17973 : 1;
	17974 : 0;
	17975 : 0;
	17976 : 0;
	17977 : 0;
	17978 : 0;
	17979 : 1;
	17980 : 1;
	17981 : 0;
	17982 : 0;
	17983 : 0;
	17984 : 0;
	17985 : 1;
	17986 : 1;
	17987 : 0;
	17988 : 0;
	17989 : 0;
	17990 : 0;
	17991 : 0;
	17992 : 1;
	17993 : 1;
	17994 : 1;
	17995 : 1;
	17996 : 1;
	17997 : 1;
	17998 : 1;
	17999 : 1;
	18000 : 1;
	18001 : 1;
	18002 : 1;
	18003 : 1;
	18004 : 1;
	18005 : 1;
	18006 : 1;
	18007 : 1;
	18008 : 1;
	18009 : 0;
	18010 : 1;
	18011 : 1;
	18012 : 1;
	18013 : 1;
	18014 : 1;
	18015 : 0;
	18016 : 0;
	18017 : 0;
	18018 : 0;
	18019 : 0;
	18020 : 0;
	18021 : 1;
	18022 : 1;
	18023 : 0;
	18024 : 0;
	18025 : 0;
	18026 : 0;
	18027 : 0;
	18028 : 0;
	18029 : 1;
	18030 : 0;
	18031 : 1;
	18032 : 1;
	18033 : 0;
	18034 : 1;
	18035 : 0;
	18036 : 1;
	18037 : 1;
	18038 : 0;
	18039 : 1;
	18040 : 1;
	18041 : 0;
	18042 : 0;
	18043 : 1;
	18044 : 1;
	18045 : 1;
	18046 : 0;
	18047 : 0;
	18048 : 1;
	18049 : 1;
	18050 : 1;
	18051 : 0;
	18052 : 1;
	18053 : 0;
	18054 : 1;
	18055 : 1;
	18056 : 1;
	18057 : 0;
	18058 : 1;
	18059 : 0;
	18060 : 1;
	18061 : 1;
	18062 : 1;
	18063 : 0;
	18064 : 1;
	18065 : 1;
	18066 : 1;
	18067 : 1;
	18068 : 1;
	18069 : 1;
	18070 : 0;
	18071 : 1;
	18072 : 1;
	18073 : 1;
	18074 : 1;
	18075 : 1;
	18076 : 0;
	18077 : 0;
	18078 : 0;
	18079 : 0;
	18080 : 0;
	18081 : 0;
	18082 : 1;
	18083 : 1;
	18084 : 1;
	18085 : 1;
	18086 : 1;
	18087 : 0;
	18088 : 1;
	18089 : 1;
	18090 : 1;
	18091 : 0;
	18092 : 1;
	18093 : 1;
	18094 : 1;
	18095 : 0;
	18096 : 0;
	18097 : 0;
	18098 : 0;
	18099 : 1;
	18100 : 0;
	18101 : 0;
	18102 : 1;
	18103 : 1;
	18104 : 1;
	18105 : 1;
	18106 : 1;
	18107 : 1;
	18108 : 0;
	18109 : 1;
	18110 : 1;
	18111 : 1;
	18112 : 0;
	18113 : 1;
	18114 : 0;
	18115 : 1;
	18116 : 1;
	18117 : 0;
	18118 : 1;
	18119 : 0;
	18120 : 1;
	18121 : 1;
	18122 : 1;
	18123 : 0;
	18124 : 0;
	18125 : 1;
	18126 : 1;
	18127 : 1;
	18128 : 0;
	18129 : 1;
	18130 : 1;
	18131 : 1;
	18132 : 0;
	18133 : 1;
	18134 : 0;
	18135 : 1;
	18136 : 1;
	18137 : 1;
	18138 : 0;
	18139 : 1;
	18140 : 0;
	18141 : 0;
	18142 : 1;
	18143 : 1;
	18144 : 0;
	18145 : 0;
	18146 : 0;
	18147 : 0;
	18148 : 0;
	18149 : 1;
	18150 : 1;
	18151 : 0;
	18152 : 0;
	18153 : 1;
	18154 : 1;
	18155 : 1;
	18156 : 0;
	18157 : 1;
	18158 : 0;
	18159 : 1;
	18160 : 1;
	18161 : 1;
	18162 : 0;
	18163 : 1;
	18164 : 0;
	18165 : 1;
	18166 : 1;
	18167 : 0;
	18168 : 1;
	18169 : 0;
	18170 : 0;
	18171 : 1;
	18172 : 1;
	18173 : 0;
	18174 : 0;
	18175 : 1;
	18176 : 1;
	18177 : 1;
	18178 : 0;
	18179 : 1;
	18180 : 0;
	18181 : 1;
	18182 : 0;
	18183 : 1;
	18184 : 0;
	18185 : 1;
	18186 : 1;
	18187 : 1;
	18188 : 0;
	18189 : 1;
	18190 : 0;
	18191 : 1;
	18192 : 1;
	18193 : 1;
	18194 : 0;
	18195 : 0;
	18196 : 1;
	18197 : 1;
	18198 : 0;
	18199 : 0;
	18200 : 1;
	18201 : 1;
	18202 : 1;
	18203 : 0;
	18204 : 1;
	18205 : 0;
	18206 : 1;
	18207 : 1;
	18208 : 1;
	18209 : 0;
	18210 : 1;
	18211 : 1;
	18212 : 0;
	18213 : 1;
	18214 : 0;
	18215 : 1;
	18216 : 1;
	18217 : 1;
	18218 : 0;
	18219 : 1;
	18220 : 0;
	18221 : 0;
	18222 : 1;
	18223 : 1;
	18224 : 0;
	18225 : 0;
	18226 : 0;
	18227 : 0;
	18228 : 1;
	18229 : 1;
	18230 : 1;
	18231 : 0;
	18232 : 1;
	18233 : 1;
	18234 : 1;
	18235 : 1;
	18236 : 1;
	18237 : 1;
	18238 : 1;
	18239 : 1;
	18240 : 1;
	18241 : 1;
	18242 : 1;
	18243 : 1;
	18244 : 1;
	18245 : 1;
	18246 : 1;
	18247 : 1;
	18248 : 1;
	18249 : 0;
	18250 : 1;
	18251 : 1;
	18252 : 1;
	18253 : 1;
	18254 : 1;
	18255 : 0;
	18256 : 1;
	18257 : 1;
	18258 : 1;
	18259 : 0;
	18260 : 0;
	18261 : 1;
	18262 : 1;
	18263 : 0;
	18264 : 0;
	18265 : 1;
	18266 : 1;
	18267 : 1;
	18268 : 0;
	18269 : 1;
	18270 : 0;
	18271 : 1;
	18272 : 1;
	18273 : 0;
	18274 : 1;
	18275 : 0;
	18276 : 1;
	18277 : 1;
	18278 : 0;
	18279 : 1;
	18280 : 1;
	18281 : 1;
	18282 : 0;
	18283 : 0;
	18284 : 0;
	18285 : 1;
	18286 : 0;
	18287 : 0;
	18288 : 1;
	18289 : 1;
	18290 : 1;
	18291 : 0;
	18292 : 1;
	18293 : 0;
	18294 : 1;
	18295 : 1;
	18296 : 1;
	18297 : 0;
	18298 : 1;
	18299 : 0;
	18300 : 1;
	18301 : 1;
	18302 : 1;
	18303 : 0;
	18304 : 1;
	18305 : 1;
	18306 : 1;
	18307 : 1;
	18308 : 1;
	18309 : 1;
	18310 : 0;
	18311 : 1;
	18312 : 1;
	18313 : 1;
	18314 : 1;
	18315 : 1;
	18316 : 0;
	18317 : 0;
	18318 : 1;
	18319 : 1;
	18320 : 1;
	18321 : 0;
	18322 : 1;
	18323 : 1;
	18324 : 1;
	18325 : 1;
	18326 : 1;
	18327 : 0;
	18328 : 1;
	18329 : 1;
	18330 : 1;
	18331 : 0;
	18332 : 1;
	18333 : 1;
	18334 : 1;
	18335 : 0;
	18336 : 0;
	18337 : 0;
	18338 : 0;
	18339 : 1;
	18340 : 0;
	18341 : 0;
	18342 : 1;
	18343 : 1;
	18344 : 1;
	18345 : 1;
	18346 : 1;
	18347 : 1;
	18348 : 0;
	18349 : 1;
	18350 : 1;
	18351 : 1;
	18352 : 0;
	18353 : 1;
	18354 : 0;
	18355 : 1;
	18356 : 1;
	18357 : 0;
	18358 : 1;
	18359 : 0;
	18360 : 1;
	18361 : 1;
	18362 : 1;
	18363 : 0;
	18364 : 0;
	18365 : 1;
	18366 : 1;
	18367 : 1;
	18368 : 0;
	18369 : 0;
	18370 : 0;
	18371 : 0;
	18372 : 0;
	18373 : 1;
	18374 : 1;
	18375 : 0;
	18376 : 1;
	18377 : 0;
	18378 : 1;
	18379 : 1;
	18380 : 0;
	18381 : 0;
	18382 : 0;
	18383 : 0;
	18384 : 0;
	18385 : 0;
	18386 : 0;
	18387 : 0;
	18388 : 1;
	18389 : 1;
	18390 : 1;
	18391 : 0;
	18392 : 0;
	18393 : 1;
	18394 : 1;
	18395 : 1;
	18396 : 0;
	18397 : 1;
	18398 : 0;
	18399 : 1;
	18400 : 1;
	18401 : 1;
	18402 : 0;
	18403 : 1;
	18404 : 0;
	18405 : 1;
	18406 : 1;
	18407 : 0;
	18408 : 1;
	18409 : 0;
	18410 : 0;
	18411 : 0;
	18412 : 0;
	18413 : 0;
	18414 : 0;
	18415 : 1;
	18416 : 1;
	18417 : 1;
	18418 : 0;
	18419 : 1;
	18420 : 0;
	18421 : 1;
	18422 : 0;
	18423 : 1;
	18424 : 0;
	18425 : 1;
	18426 : 1;
	18427 : 1;
	18428 : 0;
	18429 : 1;
	18430 : 0;
	18431 : 1;
	18432 : 1;
	18433 : 1;
	18434 : 0;
	18435 : 0;
	18436 : 1;
	18437 : 1;
	18438 : 0;
	18439 : 0;
	18440 : 1;
	18441 : 1;
	18442 : 1;
	18443 : 0;
	18444 : 1;
	18445 : 0;
	18446 : 0;
	18447 : 0;
	18448 : 0;
	18449 : 0;
	18450 : 1;
	18451 : 1;
	18452 : 0;
	18453 : 1;
	18454 : 0;
	18455 : 1;
	18456 : 1;
	18457 : 1;
	18458 : 0;
	18459 : 1;
	18460 : 0;
	18461 : 0;
	18462 : 0;
	18463 : 0;
	18464 : 0;
	18465 : 0;
	18466 : 0;
	18467 : 0;
	18468 : 1;
	18469 : 1;
	18470 : 1;
	18471 : 0;
	18472 : 1;
	18473 : 1;
	18474 : 1;
	18475 : 1;
	18476 : 1;
	18477 : 1;
	18478 : 1;
	18479 : 1;
	18480 : 1;
	18481 : 1;
	18482 : 1;
	18483 : 1;
	18484 : 1;
	18485 : 1;
	18486 : 1;
	18487 : 1;
	18488 : 1;
	18489 : 0;
	18490 : 1;
	18491 : 1;
	18492 : 1;
	18493 : 0;
	18494 : 1;
	18495 : 0;
	18496 : 1;
	18497 : 1;
	18498 : 1;
	18499 : 0;
	18500 : 0;
	18501 : 1;
	18502 : 1;
	18503 : 0;
	18504 : 0;
	18505 : 1;
	18506 : 1;
	18507 : 1;
	18508 : 0;
	18509 : 1;
	18510 : 0;
	18511 : 1;
	18512 : 1;
	18513 : 0;
	18514 : 1;
	18515 : 0;
	18516 : 1;
	18517 : 1;
	18518 : 0;
	18519 : 1;
	18520 : 1;
	18521 : 1;
	18522 : 1;
	18523 : 1;
	18524 : 0;
	18525 : 0;
	18526 : 0;
	18527 : 0;
	18528 : 1;
	18529 : 1;
	18530 : 1;
	18531 : 0;
	18532 : 1;
	18533 : 0;
	18534 : 1;
	18535 : 1;
	18536 : 1;
	18537 : 0;
	18538 : 1;
	18539 : 0;
	18540 : 1;
	18541 : 1;
	18542 : 0;
	18543 : 0;
	18544 : 1;
	18545 : 0;
	18546 : 0;
	18547 : 1;
	18548 : 1;
	18549 : 1;
	18550 : 0;
	18551 : 1;
	18552 : 1;
	18553 : 1;
	18554 : 0;
	18555 : 0;
	18556 : 0;
	18557 : 0;
	18558 : 1;
	18559 : 1;
	18560 : 1;
	18561 : 0;
	18562 : 1;
	18563 : 1;
	18564 : 1;
	18565 : 1;
	18566 : 1;
	18567 : 0;
	18568 : 1;
	18569 : 1;
	18570 : 1;
	18571 : 0;
	18572 : 1;
	18573 : 1;
	18574 : 0;
	18575 : 0;
	18576 : 0;
	18577 : 0;
	18578 : 0;
	18579 : 1;
	18580 : 0;
	18581 : 0;
	18582 : 1;
	18583 : 0;
	18584 : 0;
	18585 : 1;
	18586 : 1;
	18587 : 1;
	18588 : 0;
	18589 : 1;
	18590 : 1;
	18591 : 0;
	18592 : 0;
	18593 : 1;
	18594 : 0;
	18595 : 1;
	18596 : 1;
	18597 : 0;
	18598 : 1;
	18599 : 0;
	18600 : 1;
	18601 : 1;
	18602 : 1;
	18603 : 0;
	18604 : 0;
	18605 : 1;
	18606 : 1;
	18607 : 1;
	18608 : 0;
	18609 : 1;
	18610 : 1;
	18611 : 1;
	18612 : 1;
	18613 : 1;
	18614 : 1;
	18615 : 0;
	18616 : 1;
	18617 : 0;
	18618 : 1;
	18619 : 1;
	18620 : 0;
	18621 : 1;
	18622 : 1;
	18623 : 1;
	18624 : 1;
	18625 : 1;
	18626 : 0;
	18627 : 0;
	18628 : 1;
	18629 : 1;
	18630 : 1;
	18631 : 0;
	18632 : 0;
	18633 : 1;
	18634 : 1;
	18635 : 1;
	18636 : 0;
	18637 : 1;
	18638 : 0;
	18639 : 1;
	18640 : 1;
	18641 : 1;
	18642 : 0;
	18643 : 1;
	18644 : 0;
	18645 : 1;
	18646 : 1;
	18647 : 0;
	18648 : 1;
	18649 : 0;
	18650 : 1;
	18651 : 1;
	18652 : 1;
	18653 : 1;
	18654 : 1;
	18655 : 1;
	18656 : 1;
	18657 : 1;
	18658 : 0;
	18659 : 1;
	18660 : 0;
	18661 : 1;
	18662 : 0;
	18663 : 1;
	18664 : 0;
	18665 : 1;
	18666 : 1;
	18667 : 1;
	18668 : 0;
	18669 : 1;
	18670 : 0;
	18671 : 1;
	18672 : 1;
	18673 : 1;
	18674 : 0;
	18675 : 0;
	18676 : 1;
	18677 : 1;
	18678 : 0;
	18679 : 0;
	18680 : 1;
	18681 : 1;
	18682 : 1;
	18683 : 0;
	18684 : 1;
	18685 : 0;
	18686 : 1;
	18687 : 1;
	18688 : 1;
	18689 : 1;
	18690 : 1;
	18691 : 1;
	18692 : 0;
	18693 : 1;
	18694 : 0;
	18695 : 1;
	18696 : 1;
	18697 : 1;
	18698 : 0;
	18699 : 1;
	18700 : 0;
	18701 : 1;
	18702 : 1;
	18703 : 1;
	18704 : 1;
	18705 : 1;
	18706 : 0;
	18707 : 0;
	18708 : 1;
	18709 : 1;
	18710 : 1;
	18711 : 0;
	18712 : 1;
	18713 : 1;
	18714 : 1;
	18715 : 1;
	18716 : 1;
	18717 : 1;
	18718 : 1;
	18719 : 1;
	18720 : 1;
	18721 : 1;
	18722 : 1;
	18723 : 1;
	18724 : 1;
	18725 : 1;
	18726 : 1;
	18727 : 1;
	18728 : 1;
	18729 : 1;
	18730 : 0;
	18731 : 0;
	18732 : 0;
	18733 : 1;
	18734 : 1;
	18735 : 0;
	18736 : 1;
	18737 : 1;
	18738 : 1;
	18739 : 0;
	18740 : 0;
	18741 : 1;
	18742 : 1;
	18743 : 0;
	18744 : 0;
	18745 : 1;
	18746 : 1;
	18747 : 1;
	18748 : 0;
	18749 : 1;
	18750 : 0;
	18751 : 1;
	18752 : 1;
	18753 : 0;
	18754 : 1;
	18755 : 1;
	18756 : 0;
	18757 : 0;
	18758 : 1;
	18759 : 0;
	18760 : 1;
	18761 : 0;
	18762 : 0;
	18763 : 0;
	18764 : 0;
	18765 : 0;
	18766 : 0;
	18767 : 0;
	18768 : 1;
	18769 : 1;
	18770 : 1;
	18771 : 0;
	18772 : 1;
	18773 : 1;
	18774 : 0;
	18775 : 0;
	18776 : 0;
	18777 : 0;
	18778 : 1;
	18779 : 1;
	18780 : 0;
	18781 : 0;
	18782 : 1;
	18783 : 0;
	18784 : 1;
	18785 : 0;
	18786 : 0;
	18787 : 1;
	18788 : 1;
	18789 : 1;
	18790 : 1;
	18791 : 0;
	18792 : 0;
	18793 : 0;
	18794 : 0;
	18795 : 1;
	18796 : 0;
	18797 : 0;
	18798 : 1;
	18799 : 1;
	18800 : 1;
	18801 : 0;
	18802 : 1;
	18803 : 1;
	18804 : 1;
	18805 : 0;
	18806 : 0;
	18807 : 0;
	18808 : 0;
	18809 : 0;
	18810 : 1;
	18811 : 1;
	18812 : 0;
	18813 : 0;
	18814 : 0;
	18815 : 0;
	18816 : 0;
	18817 : 0;
	18818 : 0;
	18819 : 1;
	18820 : 0;
	18821 : 0;
	18822 : 1;
	18823 : 0;
	18824 : 0;
	18825 : 1;
	18826 : 1;
	18827 : 1;
	18828 : 1;
	18829 : 0;
	18830 : 0;
	18831 : 1;
	18832 : 0;
	18833 : 1;
	18834 : 0;
	18835 : 1;
	18836 : 1;
	18837 : 0;
	18838 : 1;
	18839 : 1;
	18840 : 0;
	18841 : 0;
	18842 : 0;
	18843 : 0;
	18844 : 0;
	18845 : 1;
	18846 : 1;
	18847 : 1;
	18848 : 1;
	18849 : 0;
	18850 : 0;
	18851 : 0;
	18852 : 0;
	18853 : 1;
	18854 : 1;
	18855 : 1;
	18856 : 0;
	18857 : 1;
	18858 : 1;
	18859 : 1;
	18860 : 1;
	18861 : 0;
	18862 : 0;
	18863 : 0;
	18864 : 0;
	18865 : 0;
	18866 : 0;
	18867 : 0;
	18868 : 1;
	18869 : 1;
	18870 : 1;
	18871 : 1;
	18872 : 0;
	18873 : 0;
	18874 : 0;
	18875 : 0;
	18876 : 0;
	18877 : 1;
	18878 : 1;
	18879 : 0;
	18880 : 0;
	18881 : 0;
	18882 : 1;
	18883 : 1;
	18884 : 0;
	18885 : 1;
	18886 : 1;
	18887 : 0;
	18888 : 1;
	18889 : 1;
	18890 : 0;
	18891 : 0;
	18892 : 0;
	18893 : 0;
	18894 : 0;
	18895 : 1;
	18896 : 1;
	18897 : 1;
	18898 : 1;
	18899 : 0;
	18900 : 1;
	18901 : 0;
	18902 : 1;
	18903 : 1;
	18904 : 0;
	18905 : 1;
	18906 : 1;
	18907 : 1;
	18908 : 0;
	18909 : 1;
	18910 : 1;
	18911 : 0;
	18912 : 0;
	18913 : 0;
	18914 : 0;
	18915 : 1;
	18916 : 1;
	18917 : 1;
	18918 : 0;
	18919 : 0;
	18920 : 1;
	18921 : 1;
	18922 : 1;
	18923 : 0;
	18924 : 1;
	18925 : 1;
	18926 : 0;
	18927 : 0;
	18928 : 0;
	18929 : 0;
	18930 : 1;
	18931 : 1;
	18932 : 0;
	18933 : 1;
	18934 : 0;
	18935 : 0;
	18936 : 0;
	18937 : 0;
	18938 : 1;
	18939 : 1;
	18940 : 1;
	18941 : 0;
	18942 : 0;
	18943 : 0;
	18944 : 0;
	18945 : 0;
	18946 : 1;
	18947 : 0;
	18948 : 0;
	18949 : 0;
	18950 : 0;
	18951 : 0;
	18952 : 1;
	18953 : 1;
	18954 : 1;
	18955 : 1;
	18956 : 1;
	18957 : 1;
	18958 : 1;
	18959 : 1;
	18960 : 1;
	18961 : 1;
	18962 : 1;
	18963 : 1;
	18964 : 1;
	18965 : 1;
	18966 : 1;
	18967 : 1;
	18968 : 1;
	18969 : 1;
	18970 : 1;
	18971 : 1;
	18972 : 1;
	18973 : 1;
	18974 : 1;
	18975 : 1;
	18976 : 1;
	18977 : 1;
	18978 : 1;
	18979 : 1;
	18980 : 1;
	18981 : 1;
	18982 : 1;
	18983 : 1;
	18984 : 1;
	18985 : 1;
	18986 : 1;
	18987 : 1;
	18988 : 1;
	18989 : 1;
	18990 : 1;
	18991 : 1;
	18992 : 1;
	18993 : 1;
	18994 : 1;
	18995 : 1;
	18996 : 1;
	18997 : 1;
	18998 : 1;
	18999 : 1;
	19000 : 1;
	19001 : 1;
	19002 : 1;
	19003 : 1;
	19004 : 1;
	19005 : 1;
	19006 : 1;
	19007 : 1;
	19008 : 1;
	19009 : 1;
	19010 : 1;
	19011 : 1;
	19012 : 1;
	19013 : 1;
	19014 : 1;
	19015 : 1;
	19016 : 1;
	19017 : 0;
	19018 : 1;
	19019 : 1;
	19020 : 1;
	19021 : 1;
	19022 : 1;
	19023 : 1;
	19024 : 1;
	19025 : 1;
	19026 : 0;
	19027 : 1;
	19028 : 1;
	19029 : 1;
	19030 : 1;
	19031 : 1;
	19032 : 1;
	19033 : 1;
	19034 : 1;
	19035 : 1;
	19036 : 1;
	19037 : 1;
	19038 : 1;
	19039 : 1;
	19040 : 1;
	19041 : 1;
	19042 : 1;
	19043 : 1;
	19044 : 1;
	19045 : 1;
	19046 : 1;
	19047 : 1;
	19048 : 1;
	19049 : 1;
	19050 : 1;
	19051 : 1;
	19052 : 1;
	19053 : 1;
	19054 : 1;
	19055 : 1;
	19056 : 1;
	19057 : 1;
	19058 : 1;
	19059 : 1;
	19060 : 1;
	19061 : 1;
	19062 : 1;
	19063 : 1;
	19064 : 0;
	19065 : 1;
	19066 : 1;
	19067 : 1;
	19068 : 1;
	19069 : 1;
	19070 : 1;
	19071 : 1;
	19072 : 1;
	19073 : 1;
	19074 : 1;
	19075 : 1;
	19076 : 1;
	19077 : 1;
	19078 : 1;
	19079 : 1;
	19080 : 1;
	19081 : 1;
	19082 : 1;
	19083 : 1;
	19084 : 1;
	19085 : 1;
	19086 : 1;
	19087 : 1;
	19088 : 1;
	19089 : 1;
	19090 : 1;
	19091 : 1;
	19092 : 1;
	19093 : 1;
	19094 : 1;
	19095 : 1;
	19096 : 1;
	19097 : 1;
	19098 : 1;
	19099 : 1;
	19100 : 1;
	19101 : 1;
	19102 : 1;
	19103 : 1;
	19104 : 1;
	19105 : 1;
	19106 : 1;
	19107 : 1;
	19108 : 1;
	19109 : 1;
	19110 : 1;
	19111 : 1;
	19112 : 1;
	19113 : 1;
	19114 : 1;
	19115 : 1;
	19116 : 0;
	19117 : 1;
	19118 : 1;
	19119 : 1;
	19120 : 1;
	19121 : 1;
	19122 : 1;
	19123 : 1;
	19124 : 1;
	19125 : 1;
	19126 : 1;
	19127 : 1;
	19128 : 1;
	19129 : 1;
	19130 : 1;
	19131 : 1;
	19132 : 1;
	19133 : 1;
	19134 : 1;
	19135 : 1;
	19136 : 1;
	19137 : 1;
	19138 : 1;
	19139 : 1;
	19140 : 1;
	19141 : 1;
	19142 : 1;
	19143 : 1;
	19144 : 1;
	19145 : 1;
	19146 : 1;
	19147 : 1;
	19148 : 1;
	19149 : 1;
	19150 : 1;
	19151 : 1;
	19152 : 1;
	19153 : 1;
	19154 : 1;
	19155 : 1;
	19156 : 1;
	19157 : 1;
	19158 : 1;
	19159 : 1;
	19160 : 1;
	19161 : 1;
	19162 : 1;
	19163 : 1;
	19164 : 1;
	19165 : 1;
	19166 : 1;
	19167 : 1;
	19168 : 1;
	19169 : 1;
	19170 : 1;
	19171 : 1;
	19172 : 1;
	19173 : 1;
	19174 : 0;
	19175 : 1;
	19176 : 1;
	19177 : 1;
	19178 : 1;
	19179 : 1;
	19180 : 1;
	19181 : 1;
	19182 : 1;
	19183 : 1;
	19184 : 1;
	19185 : 1;
	19186 : 1;
	19187 : 1;
	19188 : 1;
	19189 : 1;
	19190 : 1;
	19191 : 1;
	19192 : 1;
	19193 : 1;
	19194 : 1;
	19195 : 1;
	19196 : 1;
	19197 : 1;
	19198 : 1;
	19199 : 1;
	19200 : 1;
	19201 : 1;
	19202 : 1;
	19203 : 1;
	19204 : 1;
	19205 : 1;
	19206 : 1;
	19207 : 1;
	19208 : 1;
	19209 : 1;
	19210 : 1;
	19211 : 1;
	19212 : 1;
	19213 : 1;
	19214 : 1;
	19215 : 1;
	19216 : 1;
	19217 : 1;
	19218 : 1;
	19219 : 1;
	19220 : 1;
	19221 : 1;
	19222 : 1;
	19223 : 1;
	19224 : 1;
	19225 : 1;
	19226 : 1;
	19227 : 1;
	19228 : 1;
	19229 : 1;
	19230 : 1;
	19231 : 1;
	19232 : 1;
	19233 : 1;
	19234 : 1;
	19235 : 1;
	19236 : 1;
	19237 : 1;
	19238 : 1;
	19239 : 1;
	19240 : 1;
	19241 : 1;
	19242 : 1;
	19243 : 1;
	19244 : 1;
	19245 : 1;
	19246 : 1;
	19247 : 1;
	19248 : 1;
	19249 : 1;
	19250 : 1;
	19251 : 1;
	19252 : 1;
	19253 : 0;
	19254 : 0;
	19255 : 0;
	19256 : 0;
	19257 : 1;
	19258 : 1;
	19259 : 1;
	19260 : 1;
	19261 : 1;
	19262 : 1;
	19263 : 1;
	19264 : 1;
	19265 : 0;
	19266 : 1;
	19267 : 1;
	19268 : 1;
	19269 : 1;
	19270 : 1;
	19271 : 1;
	19272 : 1;
	19273 : 1;
	19274 : 1;
	19275 : 1;
	19276 : 1;
	19277 : 1;
	19278 : 1;
	19279 : 1;
	19280 : 1;
	19281 : 1;
	19282 : 1;
	19283 : 1;
	19284 : 1;
	19285 : 1;
	19286 : 1;
	19287 : 1;
	19288 : 1;
	19289 : 1;
	19290 : 1;
	19291 : 1;
	19292 : 1;
	19293 : 1;
	19294 : 1;
	19295 : 1;
	19296 : 1;
	19297 : 1;
	19298 : 1;
	19299 : 1;
	19300 : 1;
	19301 : 1;
	19302 : 1;
	19303 : 0;
	19304 : 1;
	19305 : 1;
	19306 : 1;
	19307 : 1;
	19308 : 1;
	19309 : 1;
	19310 : 1;
	19311 : 1;
	19312 : 1;
	19313 : 1;
	19314 : 1;
	19315 : 1;
	19316 : 1;
	19317 : 1;
	19318 : 1;
	19319 : 1;
	19320 : 1;
	19321 : 1;
	19322 : 1;
	19323 : 1;
	19324 : 1;
	19325 : 1;
	19326 : 1;
	19327 : 1;
	19328 : 1;
	19329 : 1;
	19330 : 1;
	19331 : 1;
	19332 : 1;
	19333 : 1;
	19334 : 1;
	19335 : 1;
	19336 : 1;
	19337 : 1;
	19338 : 1;
	19339 : 1;
	19340 : 1;
	19341 : 1;
	19342 : 1;
	19343 : 1;
	19344 : 1;
	19345 : 1;
	19346 : 1;
	19347 : 1;
	19348 : 1;
	19349 : 1;
	19350 : 1;
	19351 : 0;
	19352 : 0;
	19353 : 0;
	19354 : 0;
	19355 : 0;
	19356 : 1;
	19357 : 1;
	19358 : 1;
	19359 : 1;
	19360 : 1;
	19361 : 1;
	19362 : 1;
	19363 : 1;
	19364 : 1;
	19365 : 1;
	19366 : 1;
	19367 : 1;
	19368 : 1;
	19369 : 1;
	19370 : 1;
	19371 : 1;
	19372 : 1;
	19373 : 1;
	19374 : 1;
	19375 : 1;
	19376 : 1;
	19377 : 1;
	19378 : 1;
	19379 : 1;
	19380 : 1;
	19381 : 1;
	19382 : 1;
	19383 : 1;
	19384 : 1;
	19385 : 1;
	19386 : 1;
	19387 : 1;
	19388 : 1;
	19389 : 1;
	19390 : 1;
	19391 : 1;
	19392 : 1;
	19393 : 1;
	19394 : 1;
	19395 : 1;
	19396 : 1;
	19397 : 1;
	19398 : 1;
	19399 : 1;
	19400 : 1;
	19401 : 1;
	19402 : 1;
	19403 : 1;
	19404 : 1;
	19405 : 1;
	19406 : 1;
	19407 : 1;
	19408 : 1;
	19409 : 1;
	19410 : 1;
	19411 : 1;
	19412 : 1;
	19413 : 1;
	19414 : 0;
	19415 : 1;
	19416 : 1;
	19417 : 1;
	19418 : 1;
	19419 : 1;
	19420 : 1;
	19421 : 1;
	19422 : 1;
	19423 : 1;
	19424 : 1;
	19425 : 1;
	19426 : 1;
	19427 : 1;
	19428 : 1;
	19429 : 1;
	19430 : 1;
	19431 : 1;
	19432 : 1;
	19433 : 1;
	19434 : 1;
	19435 : 1;
	19436 : 1;
	19437 : 1;
	19438 : 1;
	19439 : 1;
	19440 : 1;
	19441 : 1;
	19442 : 1;
	19443 : 1;
	19444 : 1;
	19445 : 1;
	19446 : 1;
	19447 : 1;
	19448 : 1;
	19449 : 1;
	19450 : 1;
	19451 : 1;
	19452 : 1;
	19453 : 1;
	19454 : 1;
	19455 : 1;
	19456 : 1;
	19457 : 1;
	19458 : 1;
	19459 : 1;
	19460 : 1;
	19461 : 1;
	19462 : 1;
	19463 : 1;
	19464 : 1;
	19465 : 1;
	19466 : 1;
	19467 : 1;
	19468 : 1;
	19469 : 1;
	19470 : 1;
	19471 : 1;
	19472 : 1;
	19473 : 1;
	19474 : 1;
	19475 : 1;
	19476 : 1;
	19477 : 1;
	19478 : 1;
	19479 : 1;
	19480 : 1;
	19481 : 1;
	19482 : 1;
	19483 : 1;
	19484 : 1;
	19485 : 1;
	19486 : 1;
	19487 : 1;
	19488 : 1;
	19489 : 1;
	19490 : 1;
	19491 : 1;
	19492 : 1;
	19493 : 1;
	19494 : 1;
	19495 : 1;
	19496 : 1;
	19497 : 1;
	19498 : 1;
	19499 : 1;
	19500 : 1;
	19501 : 1;
	19502 : 1;
	19503 : 1;
	19504 : 1;
	19505 : 1;
	19506 : 1;
	19507 : 1;
	19508 : 1;
	19509 : 1;
	19510 : 1;
	19511 : 1;
	19512 : 1;
	19513 : 1;
	19514 : 1;
	19515 : 1;
	19516 : 1;
	19517 : 1;
	19518 : 1;
	19519 : 1;
	19520 : 1;
	19521 : 1;
	19522 : 1;
	19523 : 1;
	19524 : 1;
	19525 : 1;
	19526 : 1;
	19527 : 1;
	19528 : 1;
	19529 : 1;
	19530 : 1;
	19531 : 1;
	19532 : 1;
	19533 : 1;
	19534 : 1;
	19535 : 1;
	19536 : 1;
	19537 : 1;
	19538 : 1;
	19539 : 1;
	19540 : 1;
	19541 : 1;
	19542 : 1;
	19543 : 1;
	19544 : 1;
	19545 : 1;
	19546 : 1;
	19547 : 1;
	19548 : 1;
	19549 : 1;
	19550 : 1;
	19551 : 1;
	19552 : 1;
	19553 : 1;
	19554 : 1;
	19555 : 1;
	19556 : 1;
	19557 : 1;
	19558 : 1;
	19559 : 1;
	19560 : 1;
	19561 : 1;
	19562 : 1;
	19563 : 1;
	19564 : 1;
	19565 : 1;
	19566 : 1;
	19567 : 1;
	19568 : 1;
	19569 : 1;
	19570 : 1;
	19571 : 1;
	19572 : 1;
	19573 : 1;
	19574 : 1;
	19575 : 1;
	19576 : 1;
	19577 : 1;
	19578 : 1;
	19579 : 1;
	19580 : 1;
	19581 : 1;
	19582 : 1;
	19583 : 1;
	19584 : 1;
	19585 : 1;
	19586 : 1;
	19587 : 1;
	19588 : 1;
	19589 : 1;
	19590 : 1;
	19591 : 1;
	19592 : 1;
	19593 : 1;
	19594 : 1;
	19595 : 1;
	19596 : 1;
	19597 : 1;
	19598 : 1;
	19599 : 1;
	19600 : 1;
	19601 : 1;
	19602 : 1;
	19603 : 1;
	19604 : 1;
	19605 : 1;
	19606 : 1;
	19607 : 1;
	19608 : 1;
	19609 : 1;
	19610 : 1;
	19611 : 1;
	19612 : 1;
	19613 : 1;
	19614 : 1;
	19615 : 1;
	19616 : 1;
	19617 : 1;
	19618 : 1;
	19619 : 1;
	19620 : 1;
	19621 : 1;
	19622 : 1;
	19623 : 1;
	19624 : 1;
	19625 : 1;
	19626 : 1;
	19627 : 1;
	19628 : 1;
	19629 : 1;
	19630 : 1;
	19631 : 1;
	19632 : 1;
	19633 : 1;
	19634 : 1;
	19635 : 1;
	19636 : 1;
	19637 : 1;
	19638 : 1;
	19639 : 1;
	19640 : 1;
	19641 : 1;
	19642 : 1;
	19643 : 1;
	19644 : 1;
	19645 : 1;
	19646 : 1;
	19647 : 1;
	19648 : 1;
	19649 : 1;
	19650 : 1;
	19651 : 1;
	19652 : 1;
	19653 : 1;
	19654 : 1;
	19655 : 1;
	19656 : 1;
	19657 : 1;
	19658 : 1;
	19659 : 1;
	19660 : 1;
	19661 : 1;
	19662 : 1;
	19663 : 1;
	19664 : 1;
	19665 : 1;
	19666 : 1;
	19667 : 1;
	19668 : 1;
	19669 : 1;
	19670 : 1;
	19671 : 1;
	19672 : 1;
	19673 : 1;
	19674 : 1;
	19675 : 1;
	19676 : 1;
	19677 : 1;
	19678 : 1;
	19679 : 1;
	19680 : 1;
	19681 : 1;
	19682 : 1;
	19683 : 1;
	19684 : 1;
	19685 : 1;
	19686 : 1;
	19687 : 1;
	19688 : 1;
	19689 : 1;
	19690 : 1;
	19691 : 1;
	19692 : 1;
	19693 : 1;
	19694 : 1;
	19695 : 1;
	19696 : 1;
	19697 : 1;
	19698 : 1;
	19699 : 1;
	19700 : 1;
	19701 : 1;
	19702 : 1;
	19703 : 1;
	19704 : 1;
	19705 : 1;
	19706 : 1;
	19707 : 1;
	19708 : 1;
	19709 : 1;
	19710 : 1;
	19711 : 1;
	19712 : 1;
	19713 : 1;
	19714 : 1;
	19715 : 1;
	19716 : 1;
	19717 : 1;
	19718 : 1;
	19719 : 1;
	19720 : 1;
	19721 : 1;
	19722 : 1;
	19723 : 1;
	19724 : 1;
	19725 : 1;
	19726 : 1;
	19727 : 1;
	19728 : 1;
	19729 : 1;
	19730 : 1;
	19731 : 1;
	19732 : 1;
	19733 : 1;
	19734 : 1;
	19735 : 1;
	19736 : 1;
	19737 : 1;
	19738 : 1;
	19739 : 1;
	19740 : 1;
	19741 : 1;
	19742 : 1;
	19743 : 1;
	19744 : 1;
	19745 : 1;
	19746 : 1;
	19747 : 1;
	19748 : 1;
	19749 : 1;
	19750 : 1;
	19751 : 1;
	19752 : 1;
	19753 : 1;
	19754 : 1;
	19755 : 1;
	19756 : 1;
	19757 : 1;
	19758 : 1;
	19759 : 1;
	19760 : 1;
	19761 : 1;
	19762 : 1;
	19763 : 1;
	19764 : 1;
	19765 : 1;
	19766 : 1;
	19767 : 1;
	19768 : 1;
	19769 : 1;
	19770 : 1;
	19771 : 1;
	19772 : 1;
	19773 : 1;
	19774 : 1;
	19775 : 1;
	19776 : 1;
	19777 : 1;
	19778 : 1;
	19779 : 1;
	19780 : 1;
	19781 : 1;
	19782 : 1;
	19783 : 1;
	19784 : 1;
	19785 : 1;
	19786 : 1;
	19787 : 1;
	19788 : 1;
	19789 : 1;
	19790 : 1;
	19791 : 1;
	19792 : 1;
	19793 : 1;
	19794 : 1;
	19795 : 1;
	19796 : 1;
	19797 : 1;
	19798 : 1;
	19799 : 1;
	19800 : 1;
	19801 : 1;
	19802 : 1;
	19803 : 1;
	19804 : 1;
	19805 : 1;
	19806 : 1;
	19807 : 1;
	19808 : 1;
	19809 : 1;
	19810 : 1;
	19811 : 1;
	19812 : 1;
	19813 : 1;
	19814 : 1;
	19815 : 1;
	19816 : 1;
	19817 : 1;
	19818 : 1;
	19819 : 1;
	19820 : 1;
	19821 : 1;
	19822 : 1;
	19823 : 1;
	19824 : 1;
	19825 : 1;
	19826 : 1;
	19827 : 1;
	19828 : 1;
	19829 : 1;
	19830 : 1;
	19831 : 1;
	19832 : 1;
	19833 : 1;
	19834 : 1;
	19835 : 1;
	19836 : 1;
	19837 : 1;
	19838 : 1;
	19839 : 1;
	19840 : 1;
	19841 : 1;
	19842 : 1;
	19843 : 1;
	19844 : 1;
	19845 : 1;
	19846 : 1;
	19847 : 1;
	19848 : 1;
	19849 : 1;
	19850 : 1;
	19851 : 1;
	19852 : 1;
	19853 : 1;
	19854 : 1;
	19855 : 1;
	19856 : 1;
	19857 : 1;
	19858 : 1;
	19859 : 1;
	19860 : 1;
	19861 : 1;
	19862 : 1;
	19863 : 1;
	19864 : 1;
	19865 : 1;
	19866 : 1;
	19867 : 1;
	19868 : 1;
	19869 : 1;
	19870 : 1;
	19871 : 1;
	19872 : 1;
	19873 : 1;
	19874 : 1;
	19875 : 1;
	19876 : 1;
	19877 : 1;
	19878 : 1;
	19879 : 1;
	19880 : 1;
	19881 : 1;
	19882 : 1;
	19883 : 1;
	19884 : 1;
	19885 : 1;
	19886 : 1;
	19887 : 1;
	19888 : 1;
	19889 : 1;
	19890 : 1;
	19891 : 1;
	19892 : 1;
	19893 : 1;
	19894 : 1;
	19895 : 1;
	19896 : 1;
	19897 : 1;
	19898 : 1;
	19899 : 1;
	19900 : 1;
	19901 : 1;
	19902 : 1;
	19903 : 1;
	19904 : 1;
	19905 : 1;
	19906 : 1;
	19907 : 1;
	19908 : 1;
	19909 : 1;
	19910 : 1;
	19911 : 1;
	19912 : 1;
	19913 : 1;
	19914 : 1;
	19915 : 1;
	19916 : 1;
	19917 : 1;
	19918 : 1;
	19919 : 1;
	19920 : 1;
	19921 : 1;
	19922 : 1;
	19923 : 1;
	19924 : 1;
	19925 : 1;
	19926 : 1;
	19927 : 1;
	19928 : 1;
	19929 : 1;
	19930 : 1;
	19931 : 1;
	19932 : 1;
	19933 : 1;
	19934 : 1;
	19935 : 1;
	19936 : 1;
	19937 : 1;
	19938 : 1;
	19939 : 1;
	19940 : 1;
	19941 : 1;
	19942 : 1;
	19943 : 1;
	19944 : 1;
	19945 : 1;
	19946 : 1;
	19947 : 1;
	19948 : 1;
	19949 : 1;
	19950 : 1;
	19951 : 1;
	19952 : 1;
	19953 : 1;
	19954 : 1;
	19955 : 1;
	19956 : 1;
	19957 : 1;
	19958 : 1;
	19959 : 1;
	19960 : 1;
	19961 : 1;
	19962 : 1;
	19963 : 1;
	19964 : 1;
	19965 : 1;
	19966 : 1;
	19967 : 1;
	19968 : 1;
	19969 : 1;
	19970 : 1;
	19971 : 1;
	19972 : 1;
	19973 : 1;
	19974 : 1;
	19975 : 1;
	19976 : 1;
	19977 : 1;
	19978 : 1;
	19979 : 1;
	19980 : 1;
	19981 : 1;
	19982 : 1;
	19983 : 1;
	19984 : 1;
	19985 : 1;
	19986 : 1;
	19987 : 1;
	19988 : 1;
	19989 : 1;
	19990 : 1;
	19991 : 1;
	19992 : 1;
	19993 : 1;
	19994 : 1;
	19995 : 1;
	19996 : 1;
	19997 : 1;
	19998 : 1;
	19999 : 1;
	20000 : 1;
	20001 : 1;
	20002 : 1;
	20003 : 1;
	20004 : 1;
	20005 : 1;
	20006 : 1;
	20007 : 1;
	20008 : 1;
	20009 : 1;
	20010 : 1;
	20011 : 1;
	20012 : 1;
	20013 : 1;
	20014 : 1;
	20015 : 1;
	20016 : 1;
	20017 : 1;
	20018 : 1;
	20019 : 1;
	20020 : 1;
	20021 : 1;
	20022 : 1;
	20023 : 1;
	20024 : 1;
	20025 : 1;
	20026 : 1;
	20027 : 1;
	20028 : 1;
	20029 : 1;
	20030 : 1;
	20031 : 1;
	20032 : 1;
	20033 : 1;
	20034 : 1;
	20035 : 1;
	20036 : 1;
	20037 : 1;
	20038 : 1;
	20039 : 1;
	20040 : 1;
	20041 : 1;
	20042 : 1;
	20043 : 1;
	20044 : 1;
	20045 : 1;
	20046 : 1;
	20047 : 1;
	20048 : 1;
	20049 : 1;
	20050 : 1;
	20051 : 1;
	20052 : 1;
	20053 : 1;
	20054 : 1;
	20055 : 1;
	20056 : 1;
	20057 : 1;
	20058 : 1;
	20059 : 1;
	20060 : 1;
	20061 : 1;
	20062 : 1;
	20063 : 1;
	20064 : 1;
	20065 : 1;
	20066 : 1;
	20067 : 1;
	20068 : 1;
	20069 : 1;
	20070 : 1;
	20071 : 1;
	20072 : 1;
	20073 : 1;
	20074 : 1;
	20075 : 1;
	20076 : 1;
	20077 : 1;
	20078 : 1;
	20079 : 1;
	20080 : 1;
	20081 : 1;
	20082 : 1;
	20083 : 1;
	20084 : 1;
	20085 : 1;
	20086 : 1;
	20087 : 1;
	20088 : 1;
	20089 : 1;
	20090 : 1;
	20091 : 1;
	20092 : 1;
	20093 : 1;
	20094 : 1;
	20095 : 1;
	20096 : 1;
	20097 : 1;
	20098 : 1;
	20099 : 1;
	20100 : 1;
	20101 : 1;
	20102 : 1;
	20103 : 1;
	20104 : 1;
	20105 : 1;
	20106 : 1;
	20107 : 1;
	20108 : 1;
	20109 : 1;
	20110 : 1;
	20111 : 1;
	20112 : 1;
	20113 : 1;
	20114 : 1;
	20115 : 1;
	20116 : 1;
	20117 : 1;
	20118 : 1;
	20119 : 1;
	20120 : 1;
	20121 : 1;
	20122 : 1;
	20123 : 1;
	20124 : 1;
	20125 : 1;
	20126 : 1;
	20127 : 1;
	20128 : 1;
	20129 : 1;
	20130 : 1;
	20131 : 1;
	20132 : 1;
	20133 : 1;
	20134 : 1;
	20135 : 1;
	20136 : 1;
	20137 : 1;
	20138 : 1;
	20139 : 1;
	20140 : 1;
	20141 : 1;
	20142 : 1;
	20143 : 1;
	20144 : 1;
	20145 : 1;
	20146 : 1;
	20147 : 1;
	20148 : 1;
	20149 : 1;
	20150 : 1;
	20151 : 1;
	20152 : 1;
	20153 : 1;
	20154 : 1;
	20155 : 1;
	20156 : 1;
	20157 : 1;
	20158 : 1;
	20159 : 1;
	20160 : 1;
	20161 : 1;
	20162 : 1;
	20163 : 1;
	20164 : 1;
	20165 : 1;
	20166 : 1;
	20167 : 1;
	20168 : 1;
	20169 : 1;
	20170 : 1;
	20171 : 1;
	20172 : 1;
	20173 : 1;
	20174 : 1;
	20175 : 1;
	20176 : 1;
	20177 : 1;
	20178 : 1;
	20179 : 1;
	20180 : 1;
	20181 : 1;
	20182 : 1;
	20183 : 1;
	20184 : 1;
	20185 : 1;
	20186 : 1;
	20187 : 1;
	20188 : 1;
	20189 : 1;
	20190 : 1;
	20191 : 1;
	20192 : 1;
	20193 : 1;
	20194 : 1;
	20195 : 1;
	20196 : 1;
	20197 : 1;
	20198 : 1;
	20199 : 1;
	20200 : 1;
	20201 : 1;
	20202 : 1;
	20203 : 1;
	20204 : 1;
	20205 : 1;
	20206 : 1;
	20207 : 1;
	20208 : 1;
	20209 : 1;
	20210 : 1;
	20211 : 1;
	20212 : 1;
	20213 : 1;
	20214 : 1;
	20215 : 1;
	20216 : 1;
	20217 : 1;
	20218 : 1;
	20219 : 1;
	20220 : 1;
	20221 : 1;
	20222 : 1;
	20223 : 1;
	20224 : 1;
	20225 : 1;
	20226 : 1;
	20227 : 1;
	20228 : 1;
	20229 : 1;
	20230 : 1;
	20231 : 1;
	20232 : 1;
	20233 : 1;
	20234 : 1;
	20235 : 1;
	20236 : 1;
	20237 : 1;
	20238 : 1;
	20239 : 1;
	20240 : 1;
	20241 : 1;
	20242 : 1;
	20243 : 1;
	20244 : 1;
	20245 : 1;
	20246 : 1;
	20247 : 1;
	20248 : 1;
	20249 : 1;
	20250 : 1;
	20251 : 1;
	20252 : 1;
	20253 : 1;
	20254 : 1;
	20255 : 1;
	20256 : 1;
	20257 : 1;
	20258 : 1;
	20259 : 1;
	20260 : 1;
	20261 : 1;
	20262 : 1;
	20263 : 1;
	20264 : 1;
	20265 : 1;
	20266 : 1;
	20267 : 1;
	20268 : 1;
	20269 : 1;
	20270 : 1;
	20271 : 1;
	20272 : 1;
	20273 : 1;
	20274 : 1;
	20275 : 1;
	20276 : 1;
	20277 : 1;
	20278 : 1;
	20279 : 1;
	20280 : 1;
	20281 : 1;
	20282 : 1;
	20283 : 1;
	20284 : 1;
	20285 : 1;
	20286 : 1;
	20287 : 1;
	20288 : 1;
	20289 : 1;
	20290 : 1;
	20291 : 1;
	20292 : 1;
	20293 : 1;
	20294 : 1;
	20295 : 1;
	20296 : 1;
	20297 : 1;
	20298 : 1;
	20299 : 1;
	20300 : 1;
	20301 : 1;
	20302 : 1;
	20303 : 1;
	20304 : 1;
	20305 : 1;
	20306 : 1;
	20307 : 1;
	20308 : 1;
	20309 : 1;
	20310 : 1;
	20311 : 1;
	20312 : 1;
	20313 : 1;
	20314 : 1;
	20315 : 1;
	20316 : 1;
	20317 : 1;
	20318 : 1;
	20319 : 1;
	20320 : 1;
	20321 : 1;
	20322 : 1;
	20323 : 1;
	20324 : 1;
	20325 : 1;
	20326 : 1;
	20327 : 1;
	20328 : 1;
	20329 : 1;
	20330 : 1;
	20331 : 1;
	20332 : 1;
	20333 : 1;
	20334 : 1;
	20335 : 1;
	20336 : 1;
	20337 : 1;
	20338 : 1;
	20339 : 1;
	20340 : 1;
	20341 : 1;
	20342 : 1;
	20343 : 1;
	20344 : 1;
	20345 : 1;
	20346 : 1;
	20347 : 1;
	20348 : 1;
	20349 : 1;
	20350 : 1;
	20351 : 1;
	20352 : 1;
	20353 : 1;
	20354 : 1;
	20355 : 1;
	20356 : 1;
	20357 : 1;
	20358 : 1;
	20359 : 1;
	20360 : 1;
	20361 : 1;
	20362 : 1;
	20363 : 1;
	20364 : 1;
	20365 : 1;
	20366 : 1;
	20367 : 1;
	20368 : 1;
	20369 : 1;
	20370 : 1;
	20371 : 1;
	20372 : 1;
	20373 : 1;
	20374 : 1;
	20375 : 1;
	20376 : 1;
	20377 : 1;
	20378 : 1;
	20379 : 1;
	20380 : 1;
	20381 : 1;
	20382 : 1;
	20383 : 1;
	20384 : 1;
	20385 : 1;
	20386 : 1;
	20387 : 1;
	20388 : 1;
	20389 : 1;
	20390 : 1;
	20391 : 1;
	20392 : 1;
	20393 : 1;
	20394 : 1;
	20395 : 1;
	20396 : 1;
	20397 : 1;
	20398 : 1;
	20399 : 1;
	20400 : 1;
	20401 : 1;
	20402 : 1;
	20403 : 1;
	20404 : 1;
	20405 : 1;
	20406 : 1;
	20407 : 1;
	20408 : 1;
	20409 : 1;
	20410 : 1;
	20411 : 1;
	20412 : 1;
	20413 : 1;
	20414 : 1;
	20415 : 1;
	20416 : 1;
	20417 : 1;
	20418 : 1;
	20419 : 1;
	20420 : 1;
	20421 : 1;
	20422 : 1;
	20423 : 1;
	20424 : 1;
	20425 : 1;
	20426 : 1;
	20427 : 1;
	20428 : 1;
	20429 : 1;
	20430 : 1;
	20431 : 1;
	20432 : 1;
	20433 : 1;
	20434 : 1;
	20435 : 1;
	20436 : 1;
	20437 : 1;
	20438 : 1;
	20439 : 1;
	20440 : 1;
	20441 : 1;
	20442 : 1;
	20443 : 1;
	20444 : 1;
	20445 : 1;
	20446 : 1;
	20447 : 1;
	20448 : 1;
	20449 : 1;
	20450 : 1;
	20451 : 1;
	20452 : 1;
	20453 : 1;
	20454 : 1;
	20455 : 1;
	20456 : 1;
	20457 : 1;
	20458 : 1;
	20459 : 1;
	20460 : 1;
	20461 : 1;
	20462 : 1;
	20463 : 1;
	20464 : 1;
	20465 : 1;
	20466 : 1;
	20467 : 1;
	20468 : 1;
	20469 : 1;
	20470 : 1;
	20471 : 1;
	20472 : 1;
	20473 : 1;
	20474 : 1;
	20475 : 1;
	20476 : 1;
	20477 : 1;
	20478 : 1;
	20479 : 1;
	20480 : 1;
	20481 : 1;
	20482 : 1;
	20483 : 1;
	20484 : 1;
	20485 : 1;
	20486 : 1;
	20487 : 1;
	20488 : 1;
	20489 : 1;
	20490 : 1;
	20491 : 1;
	20492 : 1;
	20493 : 1;
	20494 : 1;
	20495 : 1;
	20496 : 1;
	20497 : 1;
	20498 : 1;
	20499 : 1;
	20500 : 1;
	20501 : 1;
	20502 : 1;
	20503 : 1;
	20504 : 1;
	20505 : 1;
	20506 : 1;
	20507 : 1;
	20508 : 1;
	20509 : 1;
	20510 : 1;
	20511 : 1;
	20512 : 1;
	20513 : 1;
	20514 : 1;
	20515 : 1;
	20516 : 1;
	20517 : 1;
	20518 : 1;
	20519 : 1;
	20520 : 1;
	20521 : 1;
	20522 : 1;
	20523 : 1;
	20524 : 1;
	20525 : 1;
	20526 : 1;
	20527 : 1;
	20528 : 1;
	20529 : 1;
	20530 : 1;
	20531 : 1;
	20532 : 1;
	20533 : 1;
	20534 : 1;
	20535 : 1;
	20536 : 1;
	20537 : 1;
	20538 : 1;
	20539 : 1;
	20540 : 1;
	20541 : 1;
	20542 : 1;
	20543 : 1;
	20544 : 1;
	20545 : 1;
	20546 : 1;
	20547 : 1;
	20548 : 1;
	20549 : 1;
	20550 : 1;
	20551 : 1;
	20552 : 1;
	20553 : 1;
	20554 : 1;
	20555 : 1;
	20556 : 1;
	20557 : 1;
	20558 : 1;
	20559 : 1;
	20560 : 1;
	20561 : 1;
	20562 : 1;
	20563 : 1;
	20564 : 1;
	20565 : 1;
	20566 : 1;
	20567 : 1;
	20568 : 1;
	20569 : 1;
	20570 : 1;
	20571 : 1;
	20572 : 1;
	20573 : 1;
	20574 : 1;
	20575 : 1;
	20576 : 1;
	20577 : 1;
	20578 : 1;
	20579 : 1;
	20580 : 1;
	20581 : 1;
	20582 : 1;
	20583 : 1;
	20584 : 1;
	20585 : 1;
	20586 : 1;
	20587 : 1;
	20588 : 1;
	20589 : 1;
	20590 : 1;
	20591 : 1;
	20592 : 1;
	20593 : 1;
	20594 : 1;
	20595 : 1;
	20596 : 1;
	20597 : 1;
	20598 : 1;
	20599 : 1;
	20600 : 1;
	20601 : 1;
	20602 : 1;
	20603 : 1;
	20604 : 1;
	20605 : 1;
	20606 : 1;
	20607 : 1;
	20608 : 1;
	20609 : 1;
	20610 : 1;
	20611 : 1;
	20612 : 1;
	20613 : 1;
	20614 : 1;
	20615 : 1;
	20616 : 1;
	20617 : 1;
	20618 : 1;
	20619 : 1;
	20620 : 1;
	20621 : 1;
	20622 : 1;
	20623 : 1;
	20624 : 1;
	20625 : 1;
	20626 : 1;
	20627 : 1;
	20628 : 1;
	20629 : 1;
	20630 : 1;
	20631 : 1;
	20632 : 1;
	20633 : 1;
	20634 : 1;
	20635 : 1;
	20636 : 1;
	20637 : 1;
	20638 : 1;
	20639 : 1;
	20640 : 1;
	20641 : 1;
	20642 : 1;
	20643 : 1;
	20644 : 1;
	20645 : 1;
	20646 : 1;
	20647 : 1;
	20648 : 1;
	20649 : 1;
	20650 : 1;
	20651 : 1;
	20652 : 1;
	20653 : 1;
	20654 : 1;
	20655 : 1;
	20656 : 1;
	20657 : 1;
	20658 : 1;
	20659 : 1;
	20660 : 1;
	20661 : 1;
	20662 : 1;
	20663 : 1;
	20664 : 1;
	20665 : 1;
	20666 : 1;
	20667 : 1;
	20668 : 1;
	20669 : 1;
	20670 : 1;
	20671 : 1;
	20672 : 1;
	20673 : 1;
	20674 : 1;
	20675 : 1;
	20676 : 1;
	20677 : 1;
	20678 : 1;
	20679 : 1;
	20680 : 1;
	20681 : 1;
	20682 : 1;
	20683 : 1;
	20684 : 1;
	20685 : 1;
	20686 : 1;
	20687 : 1;
	20688 : 1;
	20689 : 1;
	20690 : 1;
	20691 : 1;
	20692 : 1;
	20693 : 1;
	20694 : 1;
	20695 : 1;
	20696 : 1;
	20697 : 1;
	20698 : 1;
	20699 : 1;
	20700 : 1;
	20701 : 1;
	20702 : 1;
	20703 : 1;
	20704 : 1;
	20705 : 1;
	20706 : 1;
	20707 : 1;
	20708 : 1;
	20709 : 1;
	20710 : 1;
	20711 : 1;
	20712 : 1;
	20713 : 1;
	20714 : 1;
	20715 : 1;
	20716 : 1;
	20717 : 1;
	20718 : 1;
	20719 : 1;
	20720 : 1;
	20721 : 1;
	20722 : 1;
	20723 : 1;
	20724 : 1;
	20725 : 1;
	20726 : 1;
	20727 : 1;
	20728 : 1;
	20729 : 1;
	20730 : 1;
	20731 : 1;
	20732 : 1;
	20733 : 1;
	20734 : 1;
	20735 : 1;
	20736 : 1;
	20737 : 1;
	20738 : 1;
	20739 : 1;
	20740 : 1;
	20741 : 1;
	20742 : 1;
	20743 : 1;
	20744 : 1;
	20745 : 1;
	20746 : 1;
	20747 : 1;
	20748 : 1;
	20749 : 1;
	20750 : 1;
	20751 : 1;
	20752 : 1;
	20753 : 1;
	20754 : 1;
	20755 : 1;
	20756 : 1;
	20757 : 1;
	20758 : 1;
	20759 : 1;
	20760 : 1;
	20761 : 1;
	20762 : 1;
	20763 : 1;
	20764 : 1;
	20765 : 1;
	20766 : 1;
	20767 : 1;
	20768 : 1;
	20769 : 1;
	20770 : 1;
	20771 : 1;
	20772 : 1;
	20773 : 1;
	20774 : 1;
	20775 : 1;
	20776 : 1;
	20777 : 1;
	20778 : 1;
	20779 : 1;
	20780 : 1;
	20781 : 1;
	20782 : 1;
	20783 : 1;
	20784 : 1;
	20785 : 1;
	20786 : 1;
	20787 : 1;
	20788 : 1;
	20789 : 1;
	20790 : 1;
	20791 : 1;
	20792 : 1;
	20793 : 1;
	20794 : 1;
	20795 : 1;
	20796 : 1;
	20797 : 1;
	20798 : 1;
	20799 : 1;
	20800 : 1;
	20801 : 1;
	20802 : 1;
	20803 : 1;
	20804 : 1;
	20805 : 1;
	20806 : 1;
	20807 : 1;
	20808 : 1;
	20809 : 1;
	20810 : 1;
	20811 : 1;
	20812 : 1;
	20813 : 1;
	20814 : 1;
	20815 : 1;
	20816 : 1;
	20817 : 1;
	20818 : 1;
	20819 : 1;
	20820 : 1;
	20821 : 1;
	20822 : 1;
	20823 : 1;
	20824 : 1;
	20825 : 1;
	20826 : 1;
	20827 : 1;
	20828 : 1;
	20829 : 1;
	20830 : 1;
	20831 : 1;
	20832 : 1;
	20833 : 1;
	20834 : 1;
	20835 : 1;
	20836 : 1;
	20837 : 1;
	20838 : 1;
	20839 : 1;
	20840 : 1;
	20841 : 1;
	20842 : 1;
	20843 : 1;
	20844 : 1;
	20845 : 1;
	20846 : 1;
	20847 : 1;
	20848 : 1;
	20849 : 1;
	20850 : 1;
	20851 : 1;
	20852 : 1;
	20853 : 1;
	20854 : 1;
	20855 : 1;
	20856 : 1;
	20857 : 1;
	20858 : 1;
	20859 : 1;
	20860 : 1;
	20861 : 1;
	20862 : 1;
	20863 : 1;
	20864 : 1;
	20865 : 1;
	20866 : 1;
	20867 : 1;
	20868 : 1;
	20869 : 1;
	20870 : 1;
	20871 : 1;
	20872 : 1;
	20873 : 1;
	20874 : 1;
	20875 : 1;
	20876 : 1;
	20877 : 1;
	20878 : 1;
	20879 : 1;
	20880 : 1;
	20881 : 1;
	20882 : 1;
	20883 : 1;
	20884 : 1;
	20885 : 1;
	20886 : 1;
	20887 : 1;
	20888 : 1;
	20889 : 1;
	20890 : 1;
	20891 : 1;
	20892 : 1;
	20893 : 1;
	20894 : 1;
	20895 : 1;
	20896 : 1;
	20897 : 1;
	20898 : 1;
	20899 : 1;
	20900 : 1;
	20901 : 1;
	20902 : 1;
	20903 : 1;
	20904 : 1;
	20905 : 1;
	20906 : 1;
	20907 : 1;
	20908 : 1;
	20909 : 1;
	20910 : 1;
	20911 : 1;
	20912 : 1;
	20913 : 1;
	20914 : 1;
	20915 : 1;
	20916 : 1;
	20917 : 1;
	20918 : 1;
	20919 : 1;
	20920 : 1;
	20921 : 1;
	20922 : 1;
	20923 : 1;
	20924 : 1;
	20925 : 1;
	20926 : 1;
	20927 : 1;
	20928 : 1;
	20929 : 1;
	20930 : 1;
	20931 : 1;
	20932 : 1;
	20933 : 1;
	20934 : 1;
	20935 : 1;
	20936 : 1;
	20937 : 1;
	20938 : 1;
	20939 : 1;
	20940 : 1;
	20941 : 1;
	20942 : 1;
	20943 : 1;
	20944 : 1;
	20945 : 1;
	20946 : 1;
	20947 : 1;
	20948 : 1;
	20949 : 1;
	20950 : 1;
	20951 : 1;
	20952 : 1;
	20953 : 1;
	20954 : 1;
	20955 : 1;
	20956 : 1;
	20957 : 1;
	20958 : 1;
	20959 : 1;
	20960 : 1;
	20961 : 1;
	20962 : 1;
	20963 : 1;
	20964 : 1;
	20965 : 1;
	20966 : 1;
	20967 : 1;
	20968 : 1;
	20969 : 1;
	20970 : 1;
	20971 : 1;
	20972 : 1;
	20973 : 1;
	20974 : 1;
	20975 : 1;
	20976 : 1;
	20977 : 1;
	20978 : 1;
	20979 : 1;
	20980 : 1;
	20981 : 1;
	20982 : 1;
	20983 : 1;
	20984 : 1;
	20985 : 1;
	20986 : 1;
	20987 : 1;
	20988 : 1;
	20989 : 1;
	20990 : 1;
	20991 : 1;
	20992 : 1;
	20993 : 1;
	20994 : 1;
	20995 : 1;
	20996 : 1;
	20997 : 1;
	20998 : 1;
	20999 : 1;
	21000 : 1;
	21001 : 1;
	21002 : 1;
	21003 : 1;
	21004 : 1;
	21005 : 1;
	21006 : 1;
	21007 : 1;
	21008 : 1;
	21009 : 1;
	21010 : 1;
	21011 : 1;
	21012 : 1;
	21013 : 1;
	21014 : 1;
	21015 : 1;
	21016 : 1;
	21017 : 1;
	21018 : 1;
	21019 : 1;
	21020 : 1;
	21021 : 1;
	21022 : 1;
	21023 : 1;
	21024 : 1;
	21025 : 1;
	21026 : 1;
	21027 : 1;
	21028 : 1;
	21029 : 1;
	21030 : 1;
	21031 : 1;
	21032 : 1;
	21033 : 1;
	21034 : 1;
	21035 : 1;
	21036 : 1;
	21037 : 1;
	21038 : 1;
	21039 : 1;
	21040 : 1;
	21041 : 1;
	21042 : 1;
	21043 : 1;
	21044 : 1;
	21045 : 1;
	21046 : 1;
	21047 : 1;
	21048 : 1;
	21049 : 1;
	21050 : 1;
	21051 : 1;
	21052 : 1;
	21053 : 1;
	21054 : 1;
	21055 : 1;
	21056 : 1;
	21057 : 1;
	21058 : 1;
	21059 : 1;
	21060 : 1;
	21061 : 1;
	21062 : 1;
	21063 : 1;
	21064 : 1;
	21065 : 1;
	21066 : 1;
	21067 : 1;
	21068 : 1;
	21069 : 1;
	21070 : 1;
	21071 : 1;
	21072 : 1;
	21073 : 1;
	21074 : 1;
	21075 : 1;
	21076 : 1;
	21077 : 1;
	21078 : 1;
	21079 : 1;
	21080 : 1;
	21081 : 1;
	21082 : 1;
	21083 : 1;
	21084 : 1;
	21085 : 1;
	21086 : 1;
	21087 : 1;
	21088 : 1;
	21089 : 1;
	21090 : 1;
	21091 : 1;
	21092 : 1;
	21093 : 1;
	21094 : 1;
	21095 : 1;
	21096 : 1;
	21097 : 1;
	21098 : 1;
	21099 : 1;
	21100 : 1;
	21101 : 1;
	21102 : 1;
	21103 : 1;
	21104 : 1;
	21105 : 1;
	21106 : 1;
	21107 : 1;
	21108 : 1;
	21109 : 1;
	21110 : 1;
	21111 : 1;
	21112 : 1;
	21113 : 1;
	21114 : 1;
	21115 : 1;
	21116 : 1;
	21117 : 1;
	21118 : 1;
	21119 : 1;
	21120 : 1;
	21121 : 1;
	21122 : 1;
	21123 : 1;
	21124 : 1;
	21125 : 1;
	21126 : 1;
	21127 : 1;
	21128 : 1;
	21129 : 1;
	21130 : 1;
	21131 : 1;
	21132 : 1;
	21133 : 1;
	21134 : 1;
	21135 : 1;
	21136 : 1;
	21137 : 1;
	21138 : 1;
	21139 : 1;
	21140 : 1;
	21141 : 1;
	21142 : 1;
	21143 : 1;
	21144 : 1;
	21145 : 1;
	21146 : 1;
	21147 : 1;
	21148 : 1;
	21149 : 1;
	21150 : 1;
	21151 : 1;
	21152 : 1;
	21153 : 1;
	21154 : 1;
	21155 : 1;
	21156 : 1;
	21157 : 1;
	21158 : 1;
	21159 : 1;
	21160 : 1;
	21161 : 1;
	21162 : 1;
	21163 : 1;
	21164 : 1;
	21165 : 1;
	21166 : 1;
	21167 : 1;
	21168 : 1;
	21169 : 1;
	21170 : 1;
	21171 : 1;
	21172 : 1;
	21173 : 1;
	21174 : 1;
	21175 : 1;
	21176 : 1;
	21177 : 1;
	21178 : 1;
	21179 : 1;
	21180 : 1;
	21181 : 1;
	21182 : 1;
	21183 : 1;
	21184 : 1;
	21185 : 1;
	21186 : 1;
	21187 : 1;
	21188 : 1;
	21189 : 1;
	21190 : 1;
	21191 : 1;
	21192 : 1;
	21193 : 1;
	21194 : 1;
	21195 : 1;
	21196 : 1;
	21197 : 1;
	21198 : 1;
	21199 : 1;
	21200 : 1;
	21201 : 1;
	21202 : 1;
	21203 : 1;
	21204 : 1;
	21205 : 1;
	21206 : 1;
	21207 : 1;
	21208 : 1;
	21209 : 1;
	21210 : 1;
	21211 : 1;
	21212 : 1;
	21213 : 1;
	21214 : 1;
	21215 : 1;
	21216 : 1;
	21217 : 1;
	21218 : 1;
	21219 : 1;
	21220 : 1;
	21221 : 1;
	21222 : 1;
	21223 : 1;
	21224 : 1;
	21225 : 1;
	21226 : 1;
	21227 : 1;
	21228 : 1;
	21229 : 1;
	21230 : 1;
	21231 : 1;
	21232 : 1;
	21233 : 1;
	21234 : 1;
	21235 : 1;
	21236 : 1;
	21237 : 1;
	21238 : 1;
	21239 : 1;
	21240 : 1;
	21241 : 1;
	21242 : 1;
	21243 : 1;
	21244 : 1;
	21245 : 1;
	21246 : 1;
	21247 : 1;
	21248 : 1;
	21249 : 1;
	21250 : 1;
	21251 : 1;
	21252 : 1;
	21253 : 1;
	21254 : 1;
	21255 : 1;
	21256 : 1;
	21257 : 1;
	21258 : 1;
	21259 : 1;
	21260 : 1;
	21261 : 1;
	21262 : 1;
	21263 : 1;
	21264 : 1;
	21265 : 1;
	21266 : 1;
	21267 : 1;
	21268 : 1;
	21269 : 1;
	21270 : 1;
	21271 : 1;
	21272 : 1;
	21273 : 1;
	21274 : 1;
	21275 : 1;
	21276 : 1;
	21277 : 1;
	21278 : 1;
	21279 : 1;
	21280 : 1;
	21281 : 1;
	21282 : 1;
	21283 : 1;
	21284 : 1;
	21285 : 1;
	21286 : 1;
	21287 : 1;
	21288 : 1;
	21289 : 1;
	21290 : 1;
	21291 : 1;
	21292 : 1;
	21293 : 1;
	21294 : 1;
	21295 : 1;
	21296 : 1;
	21297 : 1;
	21298 : 1;
	21299 : 1;
	21300 : 1;
	21301 : 1;
	21302 : 1;
	21303 : 1;
	21304 : 1;
	21305 : 1;
	21306 : 1;
	21307 : 1;
	21308 : 1;
	21309 : 1;
	21310 : 1;
	21311 : 1;
	21312 : 1;
	21313 : 1;
	21314 : 1;
	21315 : 1;
	21316 : 1;
	21317 : 1;
	21318 : 1;
	21319 : 1;
	21320 : 1;
	21321 : 1;
	21322 : 1;
	21323 : 1;
	21324 : 1;
	21325 : 1;
	21326 : 1;
	21327 : 1;
	21328 : 1;
	21329 : 1;
	21330 : 1;
	21331 : 1;
	21332 : 1;
	21333 : 1;
	21334 : 1;
	21335 : 1;
	21336 : 1;
	21337 : 1;
	21338 : 1;
	21339 : 1;
	21340 : 1;
	21341 : 1;
	21342 : 1;
	21343 : 1;
	21344 : 1;
	21345 : 1;
	21346 : 1;
	21347 : 1;
	21348 : 1;
	21349 : 1;
	21350 : 1;
	21351 : 1;
	21352 : 1;
	21353 : 1;
	21354 : 1;
	21355 : 1;
	21356 : 1;
	21357 : 1;
	21358 : 1;
	21359 : 1;
	21360 : 1;
	21361 : 1;
	21362 : 1;
	21363 : 1;
	21364 : 1;
	21365 : 1;
	21366 : 1;
	21367 : 1;
	21368 : 1;
	21369 : 1;
	21370 : 1;
	21371 : 1;
	21372 : 1;
	21373 : 1;
	21374 : 1;
	21375 : 1;
	21376 : 1;
	21377 : 1;
	21378 : 1;
	21379 : 1;
	21380 : 1;
	21381 : 1;
	21382 : 1;
	21383 : 1;
	21384 : 1;
	21385 : 1;
	21386 : 1;
	21387 : 1;
	21388 : 1;
	21389 : 1;
	21390 : 1;
	21391 : 1;
	21392 : 1;
	21393 : 1;
	21394 : 1;
	21395 : 1;
	21396 : 1;
	21397 : 1;
	21398 : 1;
	21399 : 1;
	21400 : 1;
	21401 : 1;
	21402 : 1;
	21403 : 1;
	21404 : 1;
	21405 : 1;
	21406 : 1;
	21407 : 1;
	21408 : 1;
	21409 : 1;
	21410 : 1;
	21411 : 1;
	21412 : 1;
	21413 : 1;
	21414 : 1;
	21415 : 1;
	21416 : 1;
	21417 : 1;
	21418 : 1;
	21419 : 1;
	21420 : 1;
	21421 : 1;
	21422 : 1;
	21423 : 1;
	21424 : 1;
	21425 : 1;
	21426 : 1;
	21427 : 1;
	21428 : 1;
	21429 : 1;
	21430 : 1;
	21431 : 1;
	21432 : 1;
	21433 : 1;
	21434 : 1;
	21435 : 1;
	21436 : 1;
	21437 : 1;
	21438 : 1;
	21439 : 1;
	21440 : 1;
	21441 : 1;
	21442 : 1;
	21443 : 1;
	21444 : 1;
	21445 : 1;
	21446 : 1;
	21447 : 1;
	21448 : 1;
	21449 : 1;
	21450 : 1;
	21451 : 1;
	21452 : 1;
	21453 : 1;
	21454 : 1;
	21455 : 1;
	21456 : 1;
	21457 : 1;
	21458 : 1;
	21459 : 1;
	21460 : 1;
	21461 : 1;
	21462 : 1;
	21463 : 1;
	21464 : 1;
	21465 : 1;
	21466 : 1;
	21467 : 1;
	21468 : 1;
	21469 : 1;
	21470 : 1;
	21471 : 1;
	21472 : 1;
	21473 : 1;
	21474 : 1;
	21475 : 1;
	21476 : 1;
	21477 : 1;
	21478 : 1;
	21479 : 1;
	21480 : 1;
	21481 : 1;
	21482 : 1;
	21483 : 0;
	21484 : 0;
	21485 : 0;
	21486 : 1;
	21487 : 1;
	21488 : 1;
	21489 : 1;
	21490 : 0;
	21491 : 0;
	21492 : 1;
	21493 : 1;
	21494 : 1;
	21495 : 0;
	21496 : 0;
	21497 : 0;
	21498 : 0;
	21499 : 1;
	21500 : 1;
	21501 : 0;
	21502 : 1;
	21503 : 1;
	21504 : 1;
	21505 : 1;
	21506 : 1;
	21507 : 1;
	21508 : 1;
	21509 : 1;
	21510 : 1;
	21511 : 1;
	21512 : 1;
	21513 : 1;
	21514 : 1;
	21515 : 1;
	21516 : 1;
	21517 : 1;
	21518 : 1;
	21519 : 1;
	21520 : 1;
	21521 : 1;
	21522 : 1;
	21523 : 1;
	21524 : 1;
	21525 : 1;
	21526 : 1;
	21527 : 1;
	21528 : 1;
	21529 : 1;
	21530 : 1;
	21531 : 1;
	21532 : 1;
	21533 : 1;
	21534 : 1;
	21535 : 1;
	21536 : 1;
	21537 : 1;
	21538 : 1;
	21539 : 1;
	21540 : 1;
	21541 : 1;
	21542 : 1;
	21543 : 1;
	21544 : 1;
	21545 : 1;
	21546 : 1;
	21547 : 1;
	21548 : 1;
	21549 : 1;
	21550 : 1;
	21551 : 1;
	21552 : 1;
	21553 : 1;
	21554 : 1;
	21555 : 1;
	21556 : 1;
	21557 : 1;
	21558 : 1;
	21559 : 1;
	21560 : 1;
	21561 : 1;
	21562 : 1;
	21563 : 1;
	21564 : 1;
	21565 : 1;
	21566 : 1;
	21567 : 1;
	21568 : 1;
	21569 : 1;
	21570 : 1;
	21571 : 1;
	21572 : 1;
	21573 : 1;
	21574 : 1;
	21575 : 1;
	21576 : 1;
	21577 : 1;
	21578 : 1;
	21579 : 1;
	21580 : 1;
	21581 : 1;
	21582 : 1;
	21583 : 1;
	21584 : 1;
	21585 : 1;
	21586 : 1;
	21587 : 1;
	21588 : 1;
	21589 : 1;
	21590 : 1;
	21591 : 1;
	21592 : 1;
	21593 : 1;
	21594 : 1;
	21595 : 1;
	21596 : 1;
	21597 : 1;
	21598 : 1;
	21599 : 1;
	21600 : 1;
	21601 : 1;
	21602 : 1;
	21603 : 1;
	21604 : 1;
	21605 : 1;
	21606 : 1;
	21607 : 1;
	21608 : 1;
	21609 : 1;
	21610 : 1;
	21611 : 1;
	21612 : 1;
	21613 : 1;
	21614 : 1;
	21615 : 1;
	21616 : 1;
	21617 : 1;
	21618 : 1;
	21619 : 1;
	21620 : 1;
	21621 : 1;
	21622 : 1;
	21623 : 1;
	21624 : 1;
	21625 : 1;
	21626 : 1;
	21627 : 1;
	21628 : 1;
	21629 : 1;
	21630 : 1;
	21631 : 1;
	21632 : 1;
	21633 : 1;
	21634 : 1;
	21635 : 1;
	21636 : 1;
	21637 : 1;
	21638 : 1;
	21639 : 1;
	21640 : 1;
	21641 : 1;
	21642 : 1;
	21643 : 1;
	21644 : 1;
	21645 : 1;
	21646 : 1;
	21647 : 1;
	21648 : 1;
	21649 : 1;
	21650 : 1;
	21651 : 1;
	21652 : 1;
	21653 : 1;
	21654 : 1;
	21655 : 1;
	21656 : 1;
	21657 : 1;
	21658 : 1;
	21659 : 1;
	21660 : 1;
	21661 : 1;
	21662 : 1;
	21663 : 1;
	21664 : 1;
	21665 : 1;
	21666 : 1;
	21667 : 1;
	21668 : 1;
	21669 : 1;
	21670 : 1;
	21671 : 1;
	21672 : 1;
	21673 : 1;
	21674 : 1;
	21675 : 1;
	21676 : 1;
	21677 : 1;
	21678 : 1;
	21679 : 1;
	21680 : 1;
	21681 : 1;
	21682 : 1;
	21683 : 1;
	21684 : 1;
	21685 : 1;
	21686 : 1;
	21687 : 1;
	21688 : 1;
	21689 : 1;
	21690 : 1;
	21691 : 1;
	21692 : 1;
	21693 : 1;
	21694 : 1;
	21695 : 1;
	21696 : 1;
	21697 : 1;
	21698 : 1;
	21699 : 1;
	21700 : 1;
	21701 : 1;
	21702 : 1;
	21703 : 1;
	21704 : 1;
	21705 : 1;
	21706 : 1;
	21707 : 1;
	21708 : 1;
	21709 : 1;
	21710 : 1;
	21711 : 1;
	21712 : 1;
	21713 : 1;
	21714 : 1;
	21715 : 1;
	21716 : 1;
	21717 : 1;
	21718 : 1;
	21719 : 1;
	21720 : 1;
	21721 : 1;
	21722 : 1;
	21723 : 0;
	21724 : 0;
	21725 : 0;
	21726 : 0;
	21727 : 1;
	21728 : 1;
	21729 : 0;
	21730 : 0;
	21731 : 0;
	21732 : 0;
	21733 : 1;
	21734 : 0;
	21735 : 0;
	21736 : 0;
	21737 : 0;
	21738 : 0;
	21739 : 0;
	21740 : 1;
	21741 : 0;
	21742 : 1;
	21743 : 1;
	21744 : 1;
	21745 : 1;
	21746 : 1;
	21747 : 1;
	21748 : 1;
	21749 : 1;
	21750 : 1;
	21751 : 1;
	21752 : 1;
	21753 : 1;
	21754 : 1;
	21755 : 1;
	21756 : 1;
	21757 : 1;
	21758 : 1;
	21759 : 1;
	21760 : 1;
	21761 : 1;
	21762 : 1;
	21763 : 1;
	21764 : 1;
	21765 : 1;
	21766 : 1;
	21767 : 1;
	21768 : 1;
	21769 : 1;
	21770 : 1;
	21771 : 1;
	21772 : 1;
	21773 : 1;
	21774 : 1;
	21775 : 1;
	21776 : 1;
	21777 : 1;
	21778 : 1;
	21779 : 1;
	21780 : 1;
	21781 : 1;
	21782 : 1;
	21783 : 1;
	21784 : 1;
	21785 : 1;
	21786 : 1;
	21787 : 1;
	21788 : 1;
	21789 : 1;
	21790 : 1;
	21791 : 1;
	21792 : 1;
	21793 : 1;
	21794 : 1;
	21795 : 1;
	21796 : 1;
	21797 : 1;
	21798 : 1;
	21799 : 1;
	21800 : 1;
	21801 : 1;
	21802 : 1;
	21803 : 1;
	21804 : 1;
	21805 : 1;
	21806 : 1;
	21807 : 1;
	21808 : 1;
	21809 : 1;
	21810 : 1;
	21811 : 1;
	21812 : 1;
	21813 : 1;
	21814 : 1;
	21815 : 1;
	21816 : 1;
	21817 : 1;
	21818 : 1;
	21819 : 1;
	21820 : 1;
	21821 : 1;
	21822 : 1;
	21823 : 1;
	21824 : 1;
	21825 : 1;
	21826 : 1;
	21827 : 1;
	21828 : 1;
	21829 : 1;
	21830 : 1;
	21831 : 1;
	21832 : 1;
	21833 : 1;
	21834 : 1;
	21835 : 1;
	21836 : 1;
	21837 : 1;
	21838 : 1;
	21839 : 1;
	21840 : 1;
	21841 : 1;
	21842 : 1;
	21843 : 1;
	21844 : 1;
	21845 : 1;
	21846 : 1;
	21847 : 1;
	21848 : 1;
	21849 : 1;
	21850 : 1;
	21851 : 1;
	21852 : 1;
	21853 : 1;
	21854 : 1;
	21855 : 1;
	21856 : 1;
	21857 : 1;
	21858 : 1;
	21859 : 1;
	21860 : 1;
	21861 : 1;
	21862 : 1;
	21863 : 1;
	21864 : 1;
	21865 : 1;
	21866 : 1;
	21867 : 1;
	21868 : 1;
	21869 : 1;
	21870 : 1;
	21871 : 1;
	21872 : 1;
	21873 : 1;
	21874 : 1;
	21875 : 1;
	21876 : 1;
	21877 : 1;
	21878 : 1;
	21879 : 1;
	21880 : 1;
	21881 : 1;
	21882 : 1;
	21883 : 1;
	21884 : 1;
	21885 : 1;
	21886 : 1;
	21887 : 1;
	21888 : 1;
	21889 : 1;
	21890 : 1;
	21891 : 1;
	21892 : 1;
	21893 : 1;
	21894 : 1;
	21895 : 1;
	21896 : 1;
	21897 : 1;
	21898 : 1;
	21899 : 1;
	21900 : 1;
	21901 : 1;
	21902 : 1;
	21903 : 1;
	21904 : 1;
	21905 : 1;
	21906 : 1;
	21907 : 1;
	21908 : 1;
	21909 : 1;
	21910 : 1;
	21911 : 1;
	21912 : 1;
	21913 : 1;
	21914 : 1;
	21915 : 1;
	21916 : 1;
	21917 : 1;
	21918 : 1;
	21919 : 1;
	21920 : 1;
	21921 : 1;
	21922 : 1;
	21923 : 1;
	21924 : 1;
	21925 : 1;
	21926 : 1;
	21927 : 1;
	21928 : 1;
	21929 : 1;
	21930 : 1;
	21931 : 1;
	21932 : 1;
	21933 : 1;
	21934 : 1;
	21935 : 1;
	21936 : 1;
	21937 : 1;
	21938 : 1;
	21939 : 1;
	21940 : 1;
	21941 : 1;
	21942 : 1;
	21943 : 1;
	21944 : 1;
	21945 : 1;
	21946 : 1;
	21947 : 1;
	21948 : 1;
	21949 : 1;
	21950 : 1;
	21951 : 1;
	21952 : 1;
	21953 : 1;
	21954 : 1;
	21955 : 1;
	21956 : 1;
	21957 : 1;
	21958 : 1;
	21959 : 1;
	21960 : 1;
	21961 : 1;
	21962 : 0;
	21963 : 1;
	21964 : 1;
	21965 : 1;
	21966 : 0;
	21967 : 1;
	21968 : 0;
	21969 : 1;
	21970 : 1;
	21971 : 1;
	21972 : 0;
	21973 : 0;
	21974 : 0;
	21975 : 0;
	21976 : 1;
	21977 : 1;
	21978 : 1;
	21979 : 1;
	21980 : 1;
	21981 : 0;
	21982 : 1;
	21983 : 1;
	21984 : 1;
	21985 : 1;
	21986 : 1;
	21987 : 1;
	21988 : 1;
	21989 : 1;
	21990 : 1;
	21991 : 1;
	21992 : 1;
	21993 : 1;
	21994 : 1;
	21995 : 1;
	21996 : 1;
	21997 : 1;
	21998 : 1;
	21999 : 1;
	22000 : 1;
	22001 : 1;
	22002 : 1;
	22003 : 1;
	22004 : 1;
	22005 : 1;
	22006 : 1;
	22007 : 1;
	22008 : 1;
	22009 : 1;
	22010 : 1;
	22011 : 1;
	22012 : 1;
	22013 : 1;
	22014 : 1;
	22015 : 1;
	22016 : 1;
	22017 : 1;
	22018 : 1;
	22019 : 1;
	22020 : 1;
	22021 : 1;
	22022 : 1;
	22023 : 1;
	22024 : 1;
	22025 : 1;
	22026 : 1;
	22027 : 1;
	22028 : 1;
	22029 : 1;
	22030 : 1;
	22031 : 1;
	22032 : 1;
	22033 : 1;
	22034 : 1;
	22035 : 1;
	22036 : 1;
	22037 : 1;
	22038 : 1;
	22039 : 1;
	22040 : 1;
	22041 : 1;
	22042 : 1;
	22043 : 1;
	22044 : 1;
	22045 : 1;
	22046 : 1;
	22047 : 1;
	22048 : 1;
	22049 : 1;
	22050 : 1;
	22051 : 1;
	22052 : 1;
	22053 : 1;
	22054 : 1;
	22055 : 1;
	22056 : 1;
	22057 : 1;
	22058 : 1;
	22059 : 1;
	22060 : 1;
	22061 : 1;
	22062 : 1;
	22063 : 1;
	22064 : 1;
	22065 : 1;
	22066 : 1;
	22067 : 1;
	22068 : 1;
	22069 : 1;
	22070 : 1;
	22071 : 1;
	22072 : 1;
	22073 : 1;
	22074 : 1;
	22075 : 1;
	22076 : 1;
	22077 : 1;
	22078 : 1;
	22079 : 1;
	22080 : 1;
	22081 : 1;
	22082 : 1;
	22083 : 1;
	22084 : 1;
	22085 : 1;
	22086 : 1;
	22087 : 1;
	22088 : 1;
	22089 : 1;
	22090 : 1;
	22091 : 1;
	22092 : 1;
	22093 : 1;
	22094 : 1;
	22095 : 1;
	22096 : 1;
	22097 : 1;
	22098 : 1;
	22099 : 1;
	22100 : 1;
	22101 : 1;
	22102 : 1;
	22103 : 1;
	22104 : 1;
	22105 : 1;
	22106 : 1;
	22107 : 1;
	22108 : 1;
	22109 : 1;
	22110 : 1;
	22111 : 1;
	22112 : 1;
	22113 : 1;
	22114 : 1;
	22115 : 1;
	22116 : 1;
	22117 : 1;
	22118 : 1;
	22119 : 1;
	22120 : 1;
	22121 : 1;
	22122 : 1;
	22123 : 1;
	22124 : 1;
	22125 : 1;
	22126 : 1;
	22127 : 1;
	22128 : 1;
	22129 : 1;
	22130 : 1;
	22131 : 1;
	22132 : 1;
	22133 : 1;
	22134 : 1;
	22135 : 1;
	22136 : 1;
	22137 : 1;
	22138 : 1;
	22139 : 1;
	22140 : 1;
	22141 : 1;
	22142 : 1;
	22143 : 1;
	22144 : 1;
	22145 : 1;
	22146 : 1;
	22147 : 1;
	22148 : 1;
	22149 : 1;
	22150 : 1;
	22151 : 1;
	22152 : 1;
	22153 : 1;
	22154 : 1;
	22155 : 1;
	22156 : 1;
	22157 : 1;
	22158 : 1;
	22159 : 1;
	22160 : 1;
	22161 : 1;
	22162 : 1;
	22163 : 1;
	22164 : 1;
	22165 : 1;
	22166 : 1;
	22167 : 1;
	22168 : 1;
	22169 : 1;
	22170 : 1;
	22171 : 1;
	22172 : 1;
	22173 : 1;
	22174 : 1;
	22175 : 1;
	22176 : 1;
	22177 : 1;
	22178 : 1;
	22179 : 1;
	22180 : 1;
	22181 : 1;
	22182 : 1;
	22183 : 1;
	22184 : 1;
	22185 : 1;
	22186 : 1;
	22187 : 1;
	22188 : 1;
	22189 : 1;
	22190 : 1;
	22191 : 1;
	22192 : 1;
	22193 : 1;
	22194 : 1;
	22195 : 1;
	22196 : 1;
	22197 : 1;
	22198 : 1;
	22199 : 1;
	22200 : 1;
	22201 : 1;
	22202 : 1;
	22203 : 1;
	22204 : 1;
	22205 : 1;
	22206 : 0;
	22207 : 1;
	22208 : 0;
	22209 : 1;
	22210 : 1;
	22211 : 1;
	22212 : 0;
	22213 : 0;
	22214 : 0;
	22215 : 0;
	22216 : 1;
	22217 : 1;
	22218 : 1;
	22219 : 1;
	22220 : 1;
	22221 : 0;
	22222 : 1;
	22223 : 1;
	22224 : 1;
	22225 : 1;
	22226 : 1;
	22227 : 1;
	22228 : 1;
	22229 : 1;
	22230 : 1;
	22231 : 1;
	22232 : 1;
	22233 : 1;
	22234 : 1;
	22235 : 1;
	22236 : 1;
	22237 : 1;
	22238 : 1;
	22239 : 1;
	22240 : 1;
	22241 : 1;
	22242 : 1;
	22243 : 1;
	22244 : 1;
	22245 : 1;
	22246 : 1;
	22247 : 1;
	22248 : 1;
	22249 : 1;
	22250 : 1;
	22251 : 1;
	22252 : 1;
	22253 : 1;
	22254 : 1;
	22255 : 1;
	22256 : 1;
	22257 : 1;
	22258 : 1;
	22259 : 1;
	22260 : 1;
	22261 : 1;
	22262 : 1;
	22263 : 1;
	22264 : 1;
	22265 : 1;
	22266 : 1;
	22267 : 1;
	22268 : 1;
	22269 : 1;
	22270 : 1;
	22271 : 1;
	22272 : 1;
	22273 : 1;
	22274 : 1;
	22275 : 1;
	22276 : 1;
	22277 : 1;
	22278 : 1;
	22279 : 1;
	22280 : 1;
	22281 : 1;
	22282 : 1;
	22283 : 1;
	22284 : 1;
	22285 : 1;
	22286 : 1;
	22287 : 1;
	22288 : 1;
	22289 : 1;
	22290 : 1;
	22291 : 1;
	22292 : 1;
	22293 : 1;
	22294 : 1;
	22295 : 1;
	22296 : 1;
	22297 : 1;
	22298 : 1;
	22299 : 1;
	22300 : 1;
	22301 : 1;
	22302 : 1;
	22303 : 1;
	22304 : 1;
	22305 : 1;
	22306 : 1;
	22307 : 1;
	22308 : 1;
	22309 : 1;
	22310 : 1;
	22311 : 1;
	22312 : 1;
	22313 : 1;
	22314 : 1;
	22315 : 1;
	22316 : 1;
	22317 : 1;
	22318 : 1;
	22319 : 1;
	22320 : 1;
	22321 : 1;
	22322 : 1;
	22323 : 1;
	22324 : 1;
	22325 : 1;
	22326 : 1;
	22327 : 1;
	22328 : 1;
	22329 : 1;
	22330 : 1;
	22331 : 1;
	22332 : 1;
	22333 : 1;
	22334 : 1;
	22335 : 1;
	22336 : 1;
	22337 : 1;
	22338 : 1;
	22339 : 1;
	22340 : 1;
	22341 : 1;
	22342 : 1;
	22343 : 1;
	22344 : 1;
	22345 : 1;
	22346 : 1;
	22347 : 1;
	22348 : 1;
	22349 : 1;
	22350 : 1;
	22351 : 1;
	22352 : 1;
	22353 : 1;
	22354 : 1;
	22355 : 1;
	22356 : 1;
	22357 : 1;
	22358 : 1;
	22359 : 1;
	22360 : 1;
	22361 : 1;
	22362 : 1;
	22363 : 1;
	22364 : 1;
	22365 : 1;
	22366 : 1;
	22367 : 1;
	22368 : 1;
	22369 : 1;
	22370 : 1;
	22371 : 1;
	22372 : 1;
	22373 : 1;
	22374 : 1;
	22375 : 1;
	22376 : 1;
	22377 : 1;
	22378 : 1;
	22379 : 1;
	22380 : 1;
	22381 : 1;
	22382 : 1;
	22383 : 1;
	22384 : 1;
	22385 : 1;
	22386 : 1;
	22387 : 1;
	22388 : 1;
	22389 : 1;
	22390 : 1;
	22391 : 1;
	22392 : 1;
	22393 : 1;
	22394 : 1;
	22395 : 1;
	22396 : 1;
	22397 : 1;
	22398 : 1;
	22399 : 1;
	22400 : 1;
	22401 : 1;
	22402 : 1;
	22403 : 1;
	22404 : 1;
	22405 : 1;
	22406 : 1;
	22407 : 1;
	22408 : 1;
	22409 : 1;
	22410 : 1;
	22411 : 1;
	22412 : 1;
	22413 : 1;
	22414 : 1;
	22415 : 1;
	22416 : 1;
	22417 : 1;
	22418 : 1;
	22419 : 1;
	22420 : 1;
	22421 : 1;
	22422 : 1;
	22423 : 1;
	22424 : 1;
	22425 : 1;
	22426 : 1;
	22427 : 1;
	22428 : 1;
	22429 : 1;
	22430 : 1;
	22431 : 1;
	22432 : 1;
	22433 : 1;
	22434 : 1;
	22435 : 1;
	22436 : 1;
	22437 : 1;
	22438 : 1;
	22439 : 1;
	22440 : 1;
	22441 : 1;
	22442 : 1;
	22443 : 1;
	22444 : 1;
	22445 : 1;
	22446 : 0;
	22447 : 1;
	22448 : 0;
	22449 : 0;
	22450 : 1;
	22451 : 1;
	22452 : 0;
	22453 : 1;
	22454 : 0;
	22455 : 0;
	22456 : 1;
	22457 : 1;
	22458 : 1;
	22459 : 1;
	22460 : 1;
	22461 : 0;
	22462 : 1;
	22463 : 1;
	22464 : 1;
	22465 : 1;
	22466 : 1;
	22467 : 1;
	22468 : 1;
	22469 : 1;
	22470 : 1;
	22471 : 1;
	22472 : 1;
	22473 : 1;
	22474 : 1;
	22475 : 1;
	22476 : 1;
	22477 : 1;
	22478 : 1;
	22479 : 1;
	22480 : 1;
	22481 : 1;
	22482 : 1;
	22483 : 1;
	22484 : 1;
	22485 : 1;
	22486 : 1;
	22487 : 1;
	22488 : 1;
	22489 : 1;
	22490 : 1;
	22491 : 1;
	22492 : 1;
	22493 : 1;
	22494 : 1;
	22495 : 1;
	22496 : 1;
	22497 : 1;
	22498 : 1;
	22499 : 1;
	22500 : 1;
	22501 : 1;
	22502 : 1;
	22503 : 1;
	22504 : 1;
	22505 : 1;
	22506 : 1;
	22507 : 1;
	22508 : 1;
	22509 : 1;
	22510 : 1;
	22511 : 1;
	22512 : 1;
	22513 : 1;
	22514 : 1;
	22515 : 1;
	22516 : 1;
	22517 : 1;
	22518 : 1;
	22519 : 1;
	22520 : 1;
	22521 : 1;
	22522 : 1;
	22523 : 1;
	22524 : 1;
	22525 : 1;
	22526 : 1;
	22527 : 1;
	22528 : 1;
	22529 : 1;
	22530 : 1;
	22531 : 1;
	22532 : 1;
	22533 : 1;
	22534 : 1;
	22535 : 1;
	22536 : 1;
	22537 : 1;
	22538 : 1;
	22539 : 1;
	22540 : 1;
	22541 : 1;
	22542 : 1;
	22543 : 1;
	22544 : 1;
	22545 : 1;
	22546 : 1;
	22547 : 1;
	22548 : 1;
	22549 : 1;
	22550 : 1;
	22551 : 1;
	22552 : 1;
	22553 : 1;
	22554 : 1;
	22555 : 1;
	22556 : 1;
	22557 : 1;
	22558 : 1;
	22559 : 1;
	22560 : 1;
	22561 : 1;
	22562 : 1;
	22563 : 1;
	22564 : 1;
	22565 : 1;
	22566 : 1;
	22567 : 1;
	22568 : 1;
	22569 : 1;
	22570 : 1;
	22571 : 1;
	22572 : 1;
	22573 : 1;
	22574 : 1;
	22575 : 1;
	22576 : 1;
	22577 : 1;
	22578 : 1;
	22579 : 1;
	22580 : 1;
	22581 : 1;
	22582 : 1;
	22583 : 1;
	22584 : 1;
	22585 : 1;
	22586 : 1;
	22587 : 1;
	22588 : 1;
	22589 : 1;
	22590 : 1;
	22591 : 1;
	22592 : 1;
	22593 : 1;
	22594 : 1;
	22595 : 1;
	22596 : 1;
	22597 : 1;
	22598 : 1;
	22599 : 1;
	22600 : 1;
	22601 : 1;
	22602 : 1;
	22603 : 1;
	22604 : 1;
	22605 : 1;
	22606 : 1;
	22607 : 1;
	22608 : 1;
	22609 : 1;
	22610 : 1;
	22611 : 1;
	22612 : 1;
	22613 : 1;
	22614 : 1;
	22615 : 1;
	22616 : 1;
	22617 : 1;
	22618 : 1;
	22619 : 1;
	22620 : 1;
	22621 : 1;
	22622 : 1;
	22623 : 1;
	22624 : 1;
	22625 : 1;
	22626 : 1;
	22627 : 1;
	22628 : 1;
	22629 : 1;
	22630 : 1;
	22631 : 1;
	22632 : 1;
	22633 : 1;
	22634 : 1;
	22635 : 1;
	22636 : 1;
	22637 : 1;
	22638 : 1;
	22639 : 1;
	22640 : 1;
	22641 : 1;
	22642 : 1;
	22643 : 1;
	22644 : 1;
	22645 : 1;
	22646 : 1;
	22647 : 1;
	22648 : 1;
	22649 : 1;
	22650 : 1;
	22651 : 1;
	22652 : 1;
	22653 : 1;
	22654 : 1;
	22655 : 1;
	22656 : 1;
	22657 : 1;
	22658 : 1;
	22659 : 0;
	22660 : 1;
	22661 : 1;
	22662 : 0;
	22663 : 1;
	22664 : 1;
	22665 : 0;
	22666 : 0;
	22667 : 0;
	22668 : 0;
	22669 : 1;
	22670 : 1;
	22671 : 1;
	22672 : 0;
	22673 : 0;
	22674 : 0;
	22675 : 0;
	22676 : 0;
	22677 : 0;
	22678 : 1;
	22679 : 1;
	22680 : 1;
	22681 : 1;
	22682 : 1;
	22683 : 1;
	22684 : 0;
	22685 : 0;
	22686 : 0;
	22687 : 1;
	22688 : 1;
	22689 : 0;
	22690 : 0;
	22691 : 0;
	22692 : 0;
	22693 : 1;
	22694 : 1;
	22695 : 0;
	22696 : 0;
	22697 : 0;
	22698 : 0;
	22699 : 1;
	22700 : 1;
	22701 : 0;
	22702 : 1;
	22703 : 1;
	22704 : 1;
	22705 : 1;
	22706 : 1;
	22707 : 1;
	22708 : 1;
	22709 : 1;
	22710 : 1;
	22711 : 1;
	22712 : 1;
	22713 : 1;
	22714 : 1;
	22715 : 1;
	22716 : 1;
	22717 : 1;
	22718 : 1;
	22719 : 1;
	22720 : 1;
	22721 : 1;
	22722 : 1;
	22723 : 1;
	22724 : 1;
	22725 : 1;
	22726 : 1;
	22727 : 1;
	22728 : 1;
	22729 : 1;
	22730 : 1;
	22731 : 1;
	22732 : 1;
	22733 : 1;
	22734 : 1;
	22735 : 1;
	22736 : 1;
	22737 : 1;
	22738 : 1;
	22739 : 1;
	22740 : 1;
	22741 : 1;
	22742 : 1;
	22743 : 1;
	22744 : 1;
	22745 : 1;
	22746 : 1;
	22747 : 1;
	22748 : 1;
	22749 : 1;
	22750 : 1;
	22751 : 1;
	22752 : 1;
	22753 : 1;
	22754 : 1;
	22755 : 1;
	22756 : 1;
	22757 : 1;
	22758 : 1;
	22759 : 1;
	22760 : 1;
	22761 : 1;
	22762 : 1;
	22763 : 1;
	22764 : 1;
	22765 : 1;
	22766 : 1;
	22767 : 1;
	22768 : 1;
	22769 : 1;
	22770 : 1;
	22771 : 1;
	22772 : 1;
	22773 : 1;
	22774 : 1;
	22775 : 1;
	22776 : 1;
	22777 : 1;
	22778 : 1;
	22779 : 1;
	22780 : 1;
	22781 : 1;
	22782 : 1;
	22783 : 1;
	22784 : 1;
	22785 : 1;
	22786 : 1;
	22787 : 1;
	22788 : 1;
	22789 : 1;
	22790 : 1;
	22791 : 1;
	22792 : 1;
	22793 : 1;
	22794 : 1;
	22795 : 1;
	22796 : 1;
	22797 : 1;
	22798 : 1;
	22799 : 1;
	22800 : 1;
	22801 : 1;
	22802 : 1;
	22803 : 1;
	22804 : 1;
	22805 : 1;
	22806 : 1;
	22807 : 1;
	22808 : 1;
	22809 : 1;
	22810 : 1;
	22811 : 1;
	22812 : 1;
	22813 : 1;
	22814 : 1;
	22815 : 1;
	22816 : 1;
	22817 : 1;
	22818 : 1;
	22819 : 1;
	22820 : 1;
	22821 : 1;
	22822 : 1;
	22823 : 1;
	22824 : 1;
	22825 : 1;
	22826 : 1;
	22827 : 1;
	22828 : 1;
	22829 : 1;
	22830 : 1;
	22831 : 1;
	22832 : 1;
	22833 : 1;
	22834 : 1;
	22835 : 1;
	22836 : 1;
	22837 : 1;
	22838 : 1;
	22839 : 1;
	22840 : 1;
	22841 : 1;
	22842 : 1;
	22843 : 1;
	22844 : 1;
	22845 : 1;
	22846 : 1;
	22847 : 1;
	22848 : 1;
	22849 : 1;
	22850 : 1;
	22851 : 1;
	22852 : 1;
	22853 : 1;
	22854 : 1;
	22855 : 1;
	22856 : 1;
	22857 : 1;
	22858 : 1;
	22859 : 1;
	22860 : 1;
	22861 : 1;
	22862 : 1;
	22863 : 1;
	22864 : 1;
	22865 : 1;
	22866 : 1;
	22867 : 1;
	22868 : 1;
	22869 : 1;
	22870 : 1;
	22871 : 1;
	22872 : 1;
	22873 : 1;
	22874 : 1;
	22875 : 1;
	22876 : 1;
	22877 : 1;
	22878 : 1;
	22879 : 1;
	22880 : 1;
	22881 : 1;
	22882 : 1;
	22883 : 1;
	22884 : 1;
	22885 : 1;
	22886 : 1;
	22887 : 1;
	22888 : 1;
	22889 : 1;
	22890 : 1;
	22891 : 1;
	22892 : 1;
	22893 : 1;
	22894 : 1;
	22895 : 1;
	22896 : 1;
	22897 : 1;
	22898 : 1;
	22899 : 0;
	22900 : 1;
	22901 : 1;
	22902 : 0;
	22903 : 1;
	22904 : 1;
	22905 : 0;
	22906 : 0;
	22907 : 1;
	22908 : 1;
	22909 : 1;
	22910 : 1;
	22911 : 1;
	22912 : 0;
	22913 : 0;
	22914 : 0;
	22915 : 0;
	22916 : 1;
	22917 : 0;
	22918 : 0;
	22919 : 1;
	22920 : 1;
	22921 : 1;
	22922 : 1;
	22923 : 1;
	22924 : 1;
	22925 : 1;
	22926 : 0;
	22927 : 1;
	22928 : 0;
	22929 : 1;
	22930 : 1;
	22931 : 1;
	22932 : 0;
	22933 : 0;
	22934 : 1;
	22935 : 1;
	22936 : 1;
	22937 : 1;
	22938 : 1;
	22939 : 0;
	22940 : 1;
	22941 : 0;
	22942 : 1;
	22943 : 1;
	22944 : 1;
	22945 : 1;
	22946 : 1;
	22947 : 1;
	22948 : 1;
	22949 : 1;
	22950 : 1;
	22951 : 1;
	22952 : 1;
	22953 : 1;
	22954 : 1;
	22955 : 1;
	22956 : 1;
	22957 : 1;
	22958 : 1;
	22959 : 1;
	22960 : 1;
	22961 : 1;
	22962 : 1;
	22963 : 1;
	22964 : 1;
	22965 : 1;
	22966 : 1;
	22967 : 1;
	22968 : 1;
	22969 : 1;
	22970 : 1;
	22971 : 1;
	22972 : 1;
	22973 : 1;
	22974 : 1;
	22975 : 1;
	22976 : 1;
	22977 : 1;
	22978 : 1;
	22979 : 1;
	22980 : 1;
	22981 : 1;
	22982 : 1;
	22983 : 1;
	22984 : 1;
	22985 : 1;
	22986 : 1;
	22987 : 1;
	22988 : 1;
	22989 : 1;
	22990 : 1;
	22991 : 1;
	22992 : 1;
	22993 : 1;
	22994 : 1;
	22995 : 1;
	22996 : 1;
	22997 : 1;
	22998 : 1;
	22999 : 1;
	23000 : 1;
	23001 : 1;
	23002 : 1;
	23003 : 1;
	23004 : 1;
	23005 : 1;
	23006 : 1;
	23007 : 1;
	23008 : 1;
	23009 : 1;
	23010 : 1;
	23011 : 1;
	23012 : 1;
	23013 : 1;
	23014 : 1;
	23015 : 1;
	23016 : 1;
	23017 : 1;
	23018 : 1;
	23019 : 1;
	23020 : 1;
	23021 : 1;
	23022 : 1;
	23023 : 1;
	23024 : 1;
	23025 : 1;
	23026 : 1;
	23027 : 1;
	23028 : 1;
	23029 : 1;
	23030 : 1;
	23031 : 1;
	23032 : 1;
	23033 : 1;
	23034 : 1;
	23035 : 1;
	23036 : 1;
	23037 : 1;
	23038 : 1;
	23039 : 1;
	23040 : 1;
	23041 : 1;
	23042 : 1;
	23043 : 1;
	23044 : 1;
	23045 : 1;
	23046 : 1;
	23047 : 1;
	23048 : 1;
	23049 : 1;
	23050 : 1;
	23051 : 1;
	23052 : 1;
	23053 : 1;
	23054 : 1;
	23055 : 1;
	23056 : 1;
	23057 : 1;
	23058 : 1;
	23059 : 1;
	23060 : 1;
	23061 : 1;
	23062 : 1;
	23063 : 1;
	23064 : 1;
	23065 : 1;
	23066 : 1;
	23067 : 1;
	23068 : 1;
	23069 : 1;
	23070 : 1;
	23071 : 1;
	23072 : 1;
	23073 : 1;
	23074 : 1;
	23075 : 1;
	23076 : 1;
	23077 : 1;
	23078 : 1;
	23079 : 1;
	23080 : 1;
	23081 : 1;
	23082 : 1;
	23083 : 1;
	23084 : 1;
	23085 : 1;
	23086 : 1;
	23087 : 1;
	23088 : 1;
	23089 : 1;
	23090 : 1;
	23091 : 1;
	23092 : 1;
	23093 : 1;
	23094 : 1;
	23095 : 1;
	23096 : 1;
	23097 : 1;
	23098 : 1;
	23099 : 1;
	23100 : 1;
	23101 : 1;
	23102 : 1;
	23103 : 1;
	23104 : 1;
	23105 : 1;
	23106 : 1;
	23107 : 1;
	23108 : 1;
	23109 : 1;
	23110 : 1;
	23111 : 1;
	23112 : 1;
	23113 : 1;
	23114 : 1;
	23115 : 1;
	23116 : 1;
	23117 : 1;
	23118 : 1;
	23119 : 1;
	23120 : 1;
	23121 : 1;
	23122 : 1;
	23123 : 1;
	23124 : 1;
	23125 : 1;
	23126 : 1;
	23127 : 1;
	23128 : 1;
	23129 : 1;
	23130 : 1;
	23131 : 1;
	23132 : 1;
	23133 : 1;
	23134 : 1;
	23135 : 1;
	23136 : 1;
	23137 : 1;
	23138 : 1;
	23139 : 0;
	23140 : 1;
	23141 : 1;
	23142 : 0;
	23143 : 1;
	23144 : 1;
	23145 : 1;
	23146 : 0;
	23147 : 0;
	23148 : 0;
	23149 : 1;
	23150 : 1;
	23151 : 1;
	23152 : 0;
	23153 : 0;
	23154 : 0;
	23155 : 0;
	23156 : 1;
	23157 : 0;
	23158 : 0;
	23159 : 1;
	23160 : 1;
	23161 : 1;
	23162 : 1;
	23163 : 1;
	23164 : 1;
	23165 : 1;
	23166 : 0;
	23167 : 1;
	23168 : 0;
	23169 : 1;
	23170 : 1;
	23171 : 1;
	23172 : 0;
	23173 : 0;
	23174 : 1;
	23175 : 1;
	23176 : 1;
	23177 : 1;
	23178 : 1;
	23179 : 0;
	23180 : 1;
	23181 : 1;
	23182 : 1;
	23183 : 1;
	23184 : 1;
	23185 : 1;
	23186 : 1;
	23187 : 1;
	23188 : 1;
	23189 : 1;
	23190 : 1;
	23191 : 1;
	23192 : 1;
	23193 : 1;
	23194 : 1;
	23195 : 1;
	23196 : 1;
	23197 : 1;
	23198 : 1;
	23199 : 1;
	23200 : 1;
	23201 : 1;
	23202 : 1;
	23203 : 1;
	23204 : 1;
	23205 : 1;
	23206 : 1;
	23207 : 1;
	23208 : 1;
	23209 : 1;
	23210 : 1;
	23211 : 1;
	23212 : 1;
	23213 : 1;
	23214 : 1;
	23215 : 1;
	23216 : 1;
	23217 : 1;
	23218 : 1;
	23219 : 1;
	23220 : 1;
	23221 : 1;
	23222 : 1;
	23223 : 1;
	23224 : 1;
	23225 : 1;
	23226 : 1;
	23227 : 1;
	23228 : 1;
	23229 : 1;
	23230 : 1;
	23231 : 1;
	23232 : 1;
	23233 : 1;
	23234 : 1;
	23235 : 1;
	23236 : 1;
	23237 : 1;
	23238 : 1;
	23239 : 1;
	23240 : 1;
	23241 : 1;
	23242 : 1;
	23243 : 1;
	23244 : 1;
	23245 : 1;
	23246 : 1;
	23247 : 1;
	23248 : 1;
	23249 : 1;
	23250 : 1;
	23251 : 1;
	23252 : 1;
	23253 : 1;
	23254 : 1;
	23255 : 1;
	23256 : 1;
	23257 : 1;
	23258 : 1;
	23259 : 1;
	23260 : 1;
	23261 : 1;
	23262 : 1;
	23263 : 1;
	23264 : 1;
	23265 : 1;
	23266 : 1;
	23267 : 1;
	23268 : 1;
	23269 : 1;
	23270 : 1;
	23271 : 1;
	23272 : 1;
	23273 : 1;
	23274 : 1;
	23275 : 1;
	23276 : 1;
	23277 : 1;
	23278 : 1;
	23279 : 1;
	23280 : 1;
	23281 : 1;
	23282 : 1;
	23283 : 1;
	23284 : 1;
	23285 : 1;
	23286 : 1;
	23287 : 1;
	23288 : 1;
	23289 : 1;
	23290 : 1;
	23291 : 1;
	23292 : 1;
	23293 : 1;
	23294 : 1;
	23295 : 1;
	23296 : 1;
	23297 : 1;
	23298 : 1;
	23299 : 1;
	23300 : 1;
	23301 : 1;
	23302 : 1;
	23303 : 1;
	23304 : 1;
	23305 : 1;
	23306 : 1;
	23307 : 1;
	23308 : 1;
	23309 : 1;
	23310 : 1;
	23311 : 1;
	23312 : 1;
	23313 : 1;
	23314 : 1;
	23315 : 1;
	23316 : 1;
	23317 : 1;
	23318 : 1;
	23319 : 1;
	23320 : 1;
	23321 : 1;
	23322 : 1;
	23323 : 1;
	23324 : 1;
	23325 : 1;
	23326 : 1;
	23327 : 1;
	23328 : 1;
	23329 : 1;
	23330 : 1;
	23331 : 1;
	23332 : 1;
	23333 : 1;
	23334 : 1;
	23335 : 1;
	23336 : 1;
	23337 : 1;
	23338 : 1;
	23339 : 1;
	23340 : 1;
	23341 : 1;
	23342 : 1;
	23343 : 1;
	23344 : 1;
	23345 : 1;
	23346 : 1;
	23347 : 1;
	23348 : 1;
	23349 : 1;
	23350 : 1;
	23351 : 1;
	23352 : 1;
	23353 : 1;
	23354 : 1;
	23355 : 1;
	23356 : 1;
	23357 : 1;
	23358 : 1;
	23359 : 1;
	23360 : 1;
	23361 : 1;
	23362 : 1;
	23363 : 1;
	23364 : 1;
	23365 : 1;
	23366 : 1;
	23367 : 1;
	23368 : 1;
	23369 : 1;
	23370 : 1;
	23371 : 1;
	23372 : 1;
	23373 : 1;
	23374 : 1;
	23375 : 1;
	23376 : 1;
	23377 : 1;
	23378 : 1;
	23379 : 0;
	23380 : 1;
	23381 : 1;
	23382 : 0;
	23383 : 1;
	23384 : 1;
	23385 : 1;
	23386 : 1;
	23387 : 1;
	23388 : 0;
	23389 : 0;
	23390 : 1;
	23391 : 1;
	23392 : 0;
	23393 : 0;
	23394 : 0;
	23395 : 0;
	23396 : 1;
	23397 : 0;
	23398 : 0;
	23399 : 1;
	23400 : 1;
	23401 : 1;
	23402 : 0;
	23403 : 1;
	23404 : 1;
	23405 : 1;
	23406 : 0;
	23407 : 1;
	23408 : 0;
	23409 : 1;
	23410 : 1;
	23411 : 1;
	23412 : 0;
	23413 : 0;
	23414 : 0;
	23415 : 0;
	23416 : 1;
	23417 : 1;
	23418 : 1;
	23419 : 0;
	23420 : 1;
	23421 : 0;
	23422 : 1;
	23423 : 1;
	23424 : 1;
	23425 : 1;
	23426 : 1;
	23427 : 1;
	23428 : 1;
	23429 : 1;
	23430 : 1;
	23431 : 1;
	23432 : 1;
	23433 : 1;
	23434 : 1;
	23435 : 1;
	23436 : 1;
	23437 : 1;
	23438 : 1;
	23439 : 1;
	23440 : 1;
	23441 : 1;
	23442 : 1;
	23443 : 1;
	23444 : 1;
	23445 : 1;
	23446 : 1;
	23447 : 1;
	23448 : 1;
	23449 : 1;
	23450 : 1;
	23451 : 1;
	23452 : 1;
	23453 : 1;
	23454 : 1;
	23455 : 1;
	23456 : 1;
	23457 : 1;
	23458 : 1;
	23459 : 1;
	23460 : 1;
	23461 : 1;
	23462 : 1;
	23463 : 1;
	23464 : 1;
	23465 : 1;
	23466 : 1;
	23467 : 1;
	23468 : 1;
	23469 : 1;
	23470 : 1;
	23471 : 1;
	23472 : 1;
	23473 : 1;
	23474 : 1;
	23475 : 1;
	23476 : 1;
	23477 : 1;
	23478 : 1;
	23479 : 1;
	23480 : 1;
	23481 : 1;
	23482 : 1;
	23483 : 1;
	23484 : 1;
	23485 : 1;
	23486 : 1;
	23487 : 1;
	23488 : 1;
	23489 : 1;
	23490 : 1;
	23491 : 1;
	23492 : 1;
	23493 : 1;
	23494 : 1;
	23495 : 1;
	23496 : 1;
	23497 : 1;
	23498 : 1;
	23499 : 1;
	23500 : 1;
	23501 : 1;
	23502 : 1;
	23503 : 1;
	23504 : 1;
	23505 : 1;
	23506 : 1;
	23507 : 1;
	23508 : 1;
	23509 : 1;
	23510 : 1;
	23511 : 1;
	23512 : 1;
	23513 : 1;
	23514 : 1;
	23515 : 1;
	23516 : 1;
	23517 : 1;
	23518 : 1;
	23519 : 1;
	23520 : 1;
	23521 : 1;
	23522 : 1;
	23523 : 1;
	23524 : 1;
	23525 : 1;
	23526 : 1;
	23527 : 1;
	23528 : 1;
	23529 : 1;
	23530 : 1;
	23531 : 1;
	23532 : 1;
	23533 : 1;
	23534 : 1;
	23535 : 1;
	23536 : 1;
	23537 : 1;
	23538 : 1;
	23539 : 1;
	23540 : 1;
	23541 : 1;
	23542 : 1;
	23543 : 1;
	23544 : 1;
	23545 : 1;
	23546 : 1;
	23547 : 1;
	23548 : 1;
	23549 : 1;
	23550 : 1;
	23551 : 1;
	23552 : 1;
	23553 : 1;
	23554 : 1;
	23555 : 1;
	23556 : 1;
	23557 : 1;
	23558 : 1;
	23559 : 1;
	23560 : 1;
	23561 : 1;
	23562 : 1;
	23563 : 1;
	23564 : 1;
	23565 : 1;
	23566 : 1;
	23567 : 1;
	23568 : 1;
	23569 : 1;
	23570 : 1;
	23571 : 1;
	23572 : 1;
	23573 : 1;
	23574 : 1;
	23575 : 1;
	23576 : 1;
	23577 : 1;
	23578 : 1;
	23579 : 1;
	23580 : 1;
	23581 : 1;
	23582 : 1;
	23583 : 1;
	23584 : 1;
	23585 : 1;
	23586 : 1;
	23587 : 1;
	23588 : 1;
	23589 : 1;
	23590 : 1;
	23591 : 1;
	23592 : 1;
	23593 : 1;
	23594 : 1;
	23595 : 1;
	23596 : 1;
	23597 : 1;
	23598 : 1;
	23599 : 1;
	23600 : 1;
	23601 : 1;
	23602 : 1;
	23603 : 1;
	23604 : 1;
	23605 : 1;
	23606 : 1;
	23607 : 1;
	23608 : 1;
	23609 : 1;
	23610 : 1;
	23611 : 1;
	23612 : 1;
	23613 : 1;
	23614 : 1;
	23615 : 1;
	23616 : 1;
	23617 : 1;
	23618 : 1;
	23619 : 1;
	23620 : 0;
	23621 : 0;
	23622 : 1;
	23623 : 0;
	23624 : 1;
	23625 : 0;
	23626 : 0;
	23627 : 0;
	23628 : 0;
	23629 : 0;
	23630 : 1;
	23631 : 1;
	23632 : 0;
	23633 : 0;
	23634 : 0;
	23635 : 0;
	23636 : 1;
	23637 : 0;
	23638 : 0;
	23639 : 1;
	23640 : 1;
	23641 : 1;
	23642 : 1;
	23643 : 0;
	23644 : 0;
	23645 : 0;
	23646 : 1;
	23647 : 1;
	23648 : 1;
	23649 : 0;
	23650 : 0;
	23651 : 0;
	23652 : 0;
	23653 : 1;
	23654 : 1;
	23655 : 0;
	23656 : 0;
	23657 : 0;
	23658 : 0;
	23659 : 1;
	23660 : 1;
	23661 : 0;
	23662 : 1;
	23663 : 1;
	23664 : 1;
	23665 : 1;
	23666 : 1;
	23667 : 1;
	23668 : 1;
	23669 : 1;
	23670 : 1;
	23671 : 1;
	23672 : 1;
	23673 : 1;
	23674 : 1;
	23675 : 1;
	23676 : 1;
	23677 : 1;
	23678 : 1;
	23679 : 1;
	23680 : 1;
	23681 : 1;
	23682 : 1;
	23683 : 1;
	23684 : 1;
	23685 : 1;
	23686 : 1;
	23687 : 1;
	23688 : 1;
	23689 : 1;
	23690 : 1;
	23691 : 1;
	23692 : 1;
	23693 : 1;
	23694 : 1;
	23695 : 1;
	23696 : 1;
	23697 : 1;
	23698 : 1;
	23699 : 1;
	23700 : 1;
	23701 : 1;
	23702 : 1;
	23703 : 1;
	23704 : 1;
	23705 : 1;
	23706 : 1;
	23707 : 1;
	23708 : 1;
	23709 : 1;
	23710 : 1;
	23711 : 1;
	23712 : 1;
	23713 : 1;
	23714 : 1;
	23715 : 1;
	23716 : 1;
	23717 : 1;
	23718 : 1;
	23719 : 1;
	23720 : 1;
	23721 : 1;
	23722 : 1;
	23723 : 1;
	23724 : 1;
	23725 : 1;
	23726 : 1;
	23727 : 1;
	23728 : 1;
	23729 : 1;
	23730 : 1;
	23731 : 1;
	23732 : 1;
	23733 : 1;
	23734 : 1;
	23735 : 1;
	23736 : 1;
	23737 : 1;
	23738 : 1;
	23739 : 1;
	23740 : 1;
	23741 : 1;
	23742 : 1;
	23743 : 1;
	23744 : 1;
	23745 : 1;
	23746 : 1;
	23747 : 1;
	23748 : 1;
	23749 : 1;
	23750 : 1;
	23751 : 1;
	23752 : 1;
	23753 : 1;
	23754 : 1;
	23755 : 1;
	23756 : 1;
	23757 : 1;
	23758 : 1;
	23759 : 1;
	23760 : 1;
	23761 : 1;
	23762 : 1;
	23763 : 1;
	23764 : 1;
	23765 : 1;
	23766 : 1;
	23767 : 1;
	23768 : 1;
	23769 : 1;
	23770 : 1;
	23771 : 1;
	23772 : 1;
	23773 : 1;
	23774 : 1;
	23775 : 1;
	23776 : 1;
	23777 : 1;
	23778 : 1;
	23779 : 1;
	23780 : 1;
	23781 : 1;
	23782 : 1;
	23783 : 1;
	23784 : 1;
	23785 : 1;
	23786 : 1;
	23787 : 1;
	23788 : 1;
	23789 : 1;
	23790 : 1;
	23791 : 1;
	23792 : 1;
	23793 : 1;
	23794 : 1;
	23795 : 1;
	23796 : 1;
	23797 : 1;
	23798 : 1;
	23799 : 1;
	23800 : 1;
	23801 : 1;
	23802 : 1;
	23803 : 1;
	23804 : 1;
	23805 : 1;
	23806 : 1;
	23807 : 1;
	23808 : 1;
	23809 : 1;
	23810 : 1;
	23811 : 1;
	23812 : 1;
	23813 : 1;
	23814 : 1;
	23815 : 1;
	23816 : 1;
	23817 : 1;
	23818 : 1;
	23819 : 1;
	23820 : 1;
	23821 : 1;
	23822 : 1;
	23823 : 1;
	23824 : 1;
	23825 : 1;
	23826 : 1;
	23827 : 1;
	23828 : 1;
	23829 : 1;
	23830 : 1;
	23831 : 1;
	23832 : 1;
	23833 : 1;
	23834 : 1;
	23835 : 1;
	23836 : 1;
	23837 : 1;
	23838 : 1;
	23839 : 1;
	23840 : 1;
	23841 : 1;
	23842 : 1;
	23843 : 1;
	23844 : 1;
	23845 : 1;
	23846 : 1;
	23847 : 1;
	23848 : 1;
	23849 : 1;
	23850 : 1;
	23851 : 1;
	23852 : 1;
	23853 : 1;
	23854 : 1;
	23855 : 1;
	23856 : 1;
	23857 : 1;
	23858 : 1;
	23859 : 1;
	23860 : 1;
	23861 : 1;
	23862 : 1;
	23863 : 1;
	23864 : 1;
	23865 : 1;
	23866 : 1;
	23867 : 1;
	23868 : 1;
	23869 : 1;
	23870 : 1;
	23871 : 1;
	23872 : 1;
	23873 : 1;
	23874 : 1;
	23875 : 1;
	23876 : 1;
	23877 : 1;
	23878 : 1;
	23879 : 1;
	23880 : 1;
	23881 : 1;
	23882 : 1;
	23883 : 1;
	23884 : 1;
	23885 : 1;
	23886 : 1;
	23887 : 1;
	23888 : 1;
	23889 : 1;
	23890 : 1;
	23891 : 1;
	23892 : 1;
	23893 : 1;
	23894 : 1;
	23895 : 1;
	23896 : 1;
	23897 : 1;
	23898 : 1;
	23899 : 1;
	23900 : 1;
	23901 : 1;
	23902 : 1;
	23903 : 1;
	23904 : 1;
	23905 : 1;
	23906 : 1;
	23907 : 1;
	23908 : 1;
	23909 : 1;
	23910 : 1;
	23911 : 1;
	23912 : 1;
	23913 : 1;
	23914 : 1;
	23915 : 1;
	23916 : 1;
	23917 : 1;
	23918 : 1;
	23919 : 1;
	23920 : 1;
	23921 : 1;
	23922 : 1;
	23923 : 1;
	23924 : 1;
	23925 : 1;
	23926 : 1;
	23927 : 1;
	23928 : 1;
	23929 : 1;
	23930 : 1;
	23931 : 1;
	23932 : 1;
	23933 : 1;
	23934 : 1;
	23935 : 1;
	23936 : 1;
	23937 : 1;
	23938 : 1;
	23939 : 1;
	23940 : 1;
	23941 : 1;
	23942 : 1;
	23943 : 1;
	23944 : 1;
	23945 : 1;
	23946 : 1;
	23947 : 1;
	23948 : 1;
	23949 : 1;
	23950 : 1;
	23951 : 1;
	23952 : 1;
	23953 : 1;
	23954 : 1;
	23955 : 1;
	23956 : 1;
	23957 : 1;
	23958 : 1;
	23959 : 1;
	23960 : 1;
	23961 : 1;
	23962 : 1;
	23963 : 1;
	23964 : 1;
	23965 : 1;
	23966 : 1;
	23967 : 1;
	23968 : 1;
	23969 : 1;
	23970 : 1;
	23971 : 1;
	23972 : 1;
	23973 : 1;
	23974 : 1;
	23975 : 1;
	23976 : 1;
	23977 : 1;
	23978 : 1;
	23979 : 1;
	23980 : 1;
	23981 : 1;
	23982 : 1;
	23983 : 1;
	23984 : 1;
	23985 : 1;
	23986 : 1;
	23987 : 1;
	23988 : 1;
	23989 : 1;
	23990 : 1;
	23991 : 1;
	23992 : 1;
	23993 : 1;
	23994 : 1;
	23995 : 1;
	23996 : 1;
	23997 : 1;
	23998 : 1;
	23999 : 1;
	24000 : 1;
	24001 : 1;
	24002 : 1;
	24003 : 1;
	24004 : 1;
	24005 : 1;
	24006 : 1;
	24007 : 1;
	24008 : 1;
	24009 : 1;
	24010 : 1;
	24011 : 1;
	24012 : 1;
	24013 : 1;
	24014 : 1;
	24015 : 1;
	24016 : 1;
	24017 : 1;
	24018 : 1;
	24019 : 1;
	24020 : 1;
	24021 : 1;
	24022 : 1;
	24023 : 1;
	24024 : 1;
	24025 : 1;
	24026 : 1;
	24027 : 1;
	24028 : 1;
	24029 : 1;
	24030 : 1;
	24031 : 1;
	24032 : 1;
	24033 : 1;
	24034 : 1;
	24035 : 1;
	24036 : 1;
	24037 : 1;
	24038 : 1;
	24039 : 1;
	24040 : 1;
	24041 : 1;
	24042 : 1;
	24043 : 1;
	24044 : 1;
	24045 : 1;
	24046 : 1;
	24047 : 1;
	24048 : 1;
	24049 : 1;
	24050 : 1;
	24051 : 1;
	24052 : 1;
	24053 : 1;
	24054 : 1;
	24055 : 1;
	24056 : 1;
	24057 : 1;
	24058 : 1;
	24059 : 1;
	24060 : 1;
	24061 : 1;
	24062 : 1;
	24063 : 1;
	24064 : 1;
	24065 : 1;
	24066 : 1;
	24067 : 1;
	24068 : 1;
	24069 : 1;
	24070 : 1;
	24071 : 1;
	24072 : 1;
	24073 : 1;
	24074 : 1;
	24075 : 1;
	24076 : 1;
	24077 : 1;
	24078 : 1;
	24079 : 1;
	24080 : 1;
	24081 : 1;
	24082 : 1;
	24083 : 1;
	24084 : 1;
	24085 : 1;
	24086 : 1;
	24087 : 1;
	24088 : 1;
	24089 : 1;
	24090 : 1;
	24091 : 1;
	24092 : 1;
	24093 : 1;
	24094 : 1;
	24095 : 1;
	24096 : 1;
	24097 : 1;
	24098 : 1;
	24099 : 1;
	24100 : 1;
	24101 : 1;
	24102 : 1;
	24103 : 1;
	24104 : 1;
	24105 : 1;
	24106 : 1;
	24107 : 1;
	24108 : 1;
	24109 : 1;
	24110 : 1;
	24111 : 1;
	24112 : 1;
	24113 : 1;
	24114 : 1;
	24115 : 1;
	24116 : 1;
	24117 : 1;
	24118 : 1;
	24119 : 1;
	24120 : 1;
	24121 : 1;
	24122 : 1;
	24123 : 1;
	24124 : 1;
	24125 : 1;
	24126 : 1;
	24127 : 1;
	24128 : 1;
	24129 : 1;
	24130 : 1;
	24131 : 1;
	24132 : 1;
	24133 : 1;
	24134 : 1;
	24135 : 1;
	24136 : 1;
	24137 : 1;
	24138 : 1;
	24139 : 1;
	24140 : 1;
	24141 : 1;
	24142 : 1;
	24143 : 1;
	24144 : 1;
	24145 : 1;
	24146 : 1;
	24147 : 1;
	24148 : 1;
	24149 : 1;
	24150 : 1;
	24151 : 1;
	24152 : 1;
	24153 : 1;
	24154 : 1;
	24155 : 1;
	24156 : 1;
	24157 : 1;
	24158 : 1;
	24159 : 1;
	24160 : 1;
	24161 : 1;
	24162 : 1;
	24163 : 1;
	24164 : 1;
	24165 : 1;
	24166 : 1;
	24167 : 1;
	24168 : 1;
	24169 : 1;
	24170 : 1;
	24171 : 1;
	24172 : 1;
	24173 : 1;
	24174 : 1;
	24175 : 1;
	24176 : 1;
	24177 : 1;
	24178 : 1;
	24179 : 1;
	24180 : 1;
	24181 : 1;
	24182 : 1;
	24183 : 1;
	24184 : 1;
	24185 : 1;
	24186 : 1;
	24187 : 1;
	24188 : 1;
	24189 : 1;
	24190 : 1;
	24191 : 1;
	24192 : 1;
	24193 : 1;
	24194 : 1;
	24195 : 1;
	24196 : 1;
	24197 : 1;
	24198 : 1;
	24199 : 1;
	24200 : 1;
	24201 : 1;
	24202 : 1;
	24203 : 1;
	24204 : 1;
	24205 : 1;
	24206 : 1;
	24207 : 1;
	24208 : 1;
	24209 : 1;
	24210 : 1;
	24211 : 1;
	24212 : 1;
	24213 : 1;
	24214 : 1;
	24215 : 1;
	24216 : 1;
	24217 : 1;
	24218 : 1;
	24219 : 1;
	24220 : 1;
	24221 : 1;
	24222 : 1;
	24223 : 1;
	24224 : 1;
	24225 : 1;
	24226 : 1;
	24227 : 1;
	24228 : 1;
	24229 : 1;
	24230 : 1;
	24231 : 1;
	24232 : 1;
	24233 : 1;
	24234 : 1;
	24235 : 1;
	24236 : 1;
	24237 : 1;
	24238 : 1;
	24239 : 1;
	24240 : 1;
	24241 : 1;
	24242 : 1;
	24243 : 1;
	24244 : 1;
	24245 : 1;
	24246 : 1;
	24247 : 1;
	24248 : 1;
	24249 : 1;
	24250 : 1;
	24251 : 1;
	24252 : 1;
	24253 : 1;
	24254 : 1;
	24255 : 1;
	24256 : 1;
	24257 : 1;
	24258 : 1;
	24259 : 1;
	24260 : 1;
	24261 : 1;
	24262 : 1;
	24263 : 1;
	24264 : 1;
	24265 : 1;
	24266 : 1;
	24267 : 1;
	24268 : 1;
	24269 : 1;
	24270 : 1;
	24271 : 1;
	24272 : 1;
	24273 : 1;
	24274 : 1;
	24275 : 1;
	24276 : 1;
	24277 : 1;
	24278 : 1;
	24279 : 1;
	24280 : 1;
	24281 : 1;
	24282 : 1;
	24283 : 1;
	24284 : 1;
	24285 : 1;
	24286 : 1;
	24287 : 1;
	24288 : 1;
	24289 : 1;
	24290 : 1;
	24291 : 1;
	24292 : 1;
	24293 : 1;
	24294 : 1;
	24295 : 1;
	24296 : 1;
	24297 : 1;
	24298 : 1;
	24299 : 1;
	24300 : 1;
	24301 : 1;
	24302 : 1;
	24303 : 1;
	24304 : 1;
	24305 : 1;
	24306 : 1;
	24307 : 1;
	24308 : 1;
	24309 : 1;
	24310 : 1;
	24311 : 1;
	24312 : 1;
	24313 : 1;
	24314 : 1;
	24315 : 1;
	24316 : 1;
	24317 : 1;
	24318 : 1;
	24319 : 1;
	24320 : 1;
	24321 : 1;
	24322 : 1;
	24323 : 1;
	24324 : 1;
	24325 : 1;
	24326 : 1;
	24327 : 1;
	24328 : 1;
	24329 : 1;
	24330 : 1;
	24331 : 1;
	24332 : 1;
	24333 : 1;
	24334 : 1;
	24335 : 1;
	24336 : 1;
	24337 : 1;
	24338 : 1;
	24339 : 1;
	24340 : 1;
	24341 : 1;
	24342 : 1;
	24343 : 1;
	24344 : 1;
	24345 : 1;
	24346 : 1;
	24347 : 1;
	24348 : 1;
	24349 : 1;
	24350 : 1;
	24351 : 1;
	24352 : 1;
	24353 : 1;
	24354 : 1;
	24355 : 1;
	24356 : 1;
	24357 : 1;
	24358 : 1;
	24359 : 1;
	24360 : 1;
	24361 : 1;
	24362 : 1;
	24363 : 1;
	24364 : 1;
	24365 : 1;
	24366 : 1;
	24367 : 1;
	24368 : 1;
	24369 : 1;
	24370 : 1;
	24371 : 1;
	24372 : 1;
	24373 : 1;
	24374 : 1;
	24375 : 1;
	24376 : 1;
	24377 : 1;
	24378 : 1;
	24379 : 1;
	24380 : 1;
	24381 : 1;
	24382 : 1;
	24383 : 1;
	24384 : 1;
	24385 : 1;
	24386 : 1;
	24387 : 1;
	24388 : 1;
	24389 : 1;
	24390 : 1;
	24391 : 1;
	24392 : 1;
	24393 : 1;
	24394 : 1;
	24395 : 1;
	24396 : 1;
	24397 : 1;
	24398 : 1;
	24399 : 1;
	24400 : 1;
	24401 : 1;
	24402 : 1;
	24403 : 1;
	24404 : 1;
	24405 : 1;
	24406 : 1;
	24407 : 1;
	24408 : 1;
	24409 : 1;
	24410 : 1;
	24411 : 1;
	24412 : 1;
	24413 : 1;
	24414 : 1;
	24415 : 1;
	24416 : 1;
	24417 : 1;
	24418 : 1;
	24419 : 1;
	24420 : 1;
	24421 : 1;
	24422 : 1;
	24423 : 1;
	24424 : 1;
	24425 : 1;
	24426 : 1;
	24427 : 1;
	24428 : 1;
	24429 : 1;
	24430 : 1;
	24431 : 1;
	24432 : 1;
	24433 : 1;
	24434 : 1;
	24435 : 1;
	24436 : 1;
	24437 : 1;
	24438 : 1;
	24439 : 1;
	24440 : 1;
	24441 : 1;
	24442 : 1;
	24443 : 1;
	24444 : 1;
	24445 : 1;
	24446 : 1;
	24447 : 1;
	24448 : 1;
	24449 : 1;
	24450 : 1;
	24451 : 1;
	24452 : 1;
	24453 : 1;
	24454 : 1;
	24455 : 1;
	24456 : 1;
	24457 : 1;
	24458 : 1;
	24459 : 1;
	24460 : 1;
	24461 : 1;
	24462 : 1;
	24463 : 1;
	24464 : 1;
	24465 : 1;
	24466 : 1;
	24467 : 1;
	24468 : 1;
	24469 : 1;
	24470 : 1;
	24471 : 1;
	24472 : 1;
	24473 : 1;
	24474 : 1;
	24475 : 1;
	24476 : 1;
	24477 : 1;
	24478 : 1;
	24479 : 1;
	24480 : 1;
	24481 : 1;
	24482 : 1;
	24483 : 1;
	24484 : 1;
	24485 : 1;
	24486 : 1;
	24487 : 1;
	24488 : 1;
	24489 : 1;
	24490 : 1;
	24491 : 1;
	24492 : 1;
	24493 : 1;
	24494 : 1;
	24495 : 1;
	24496 : 1;
	24497 : 1;
	24498 : 1;
	24499 : 1;
	24500 : 1;
	24501 : 1;
	24502 : 1;
	24503 : 1;
	24504 : 1;
	24505 : 1;
	24506 : 1;
	24507 : 1;
	24508 : 1;
	24509 : 1;
	24510 : 1;
	24511 : 1;
	24512 : 1;
	24513 : 1;
	24514 : 1;
	24515 : 1;
	24516 : 1;
	24517 : 1;
	24518 : 1;
	24519 : 1;
	24520 : 1;
	24521 : 1;
	24522 : 1;
	24523 : 1;
	24524 : 1;
	24525 : 1;
	24526 : 1;
	24527 : 1;
	24528 : 1;
	24529 : 1;
	24530 : 1;
	24531 : 1;
	24532 : 1;
	24533 : 1;
	24534 : 1;
	24535 : 1;
	24536 : 1;
	24537 : 1;
	24538 : 1;
	24539 : 1;
	24540 : 1;
	24541 : 1;
	24542 : 1;
	24543 : 1;
	24544 : 1;
	24545 : 1;
	24546 : 1;
	24547 : 1;
	24548 : 1;
	24549 : 1;
	24550 : 1;
	24551 : 1;
	24552 : 1;
	24553 : 1;
	24554 : 1;
	24555 : 1;
	24556 : 1;
	24557 : 1;
	24558 : 1;
	24559 : 1;
	24560 : 1;
	24561 : 1;
	24562 : 1;
	24563 : 1;
	24564 : 1;
	24565 : 1;
	24566 : 1;
	24567 : 1;
	24568 : 1;
	24569 : 1;
	24570 : 1;
	24571 : 1;
	24572 : 1;
	24573 : 1;
	24574 : 1;
	24575 : 1;
	24576 : 1;
	24577 : 1;
	24578 : 1;
	24579 : 1;
	24580 : 1;
	24581 : 1;
	24582 : 1;
	24583 : 1;
	24584 : 1;
	24585 : 1;
	24586 : 1;
	24587 : 1;
	24588 : 1;
	24589 : 1;
	24590 : 1;
	24591 : 1;
	24592 : 1;
	24593 : 1;
	24594 : 1;
	24595 : 1;
	24596 : 1;
	24597 : 1;
	24598 : 1;
	24599 : 1;
	24600 : 1;
	24601 : 1;
	24602 : 1;
	24603 : 1;
	24604 : 1;
	24605 : 1;
	24606 : 1;
	24607 : 1;
	24608 : 1;
	24609 : 1;
	24610 : 1;
	24611 : 1;
	24612 : 1;
	24613 : 1;
	24614 : 1;
	24615 : 1;
	24616 : 1;
	24617 : 1;
	24618 : 1;
	24619 : 1;
	24620 : 1;
	24621 : 1;
	24622 : 1;
	24623 : 1;
	24624 : 1;
	24625 : 1;
	24626 : 1;
	24627 : 1;
	24628 : 1;
	24629 : 1;
	24630 : 1;
	24631 : 1;
	24632 : 1;
	24633 : 1;
	24634 : 1;
	24635 : 1;
	24636 : 1;
	24637 : 1;
	24638 : 1;
	24639 : 1;
	24640 : 1;
	24641 : 1;
	24642 : 1;
	24643 : 1;
	24644 : 1;
	24645 : 1;
	24646 : 1;
	24647 : 1;
	24648 : 1;
	24649 : 1;
	24650 : 1;
	24651 : 1;
	24652 : 1;
	24653 : 1;
	24654 : 1;
	24655 : 1;
	24656 : 1;
	24657 : 1;
	24658 : 1;
	24659 : 1;
	24660 : 1;
	24661 : 1;
	24662 : 1;
	24663 : 1;
	24664 : 1;
	24665 : 1;
	24666 : 1;
	24667 : 1;
	24668 : 1;
	24669 : 1;
	24670 : 1;
	24671 : 1;
	24672 : 1;
	24673 : 1;
	24674 : 1;
	24675 : 1;
	24676 : 1;
	24677 : 1;
	24678 : 1;
	24679 : 1;
	24680 : 1;
	24681 : 1;
	24682 : 1;
	24683 : 1;
	24684 : 1;
	24685 : 1;
	24686 : 1;
	24687 : 1;
	24688 : 1;
	24689 : 1;
	24690 : 1;
	24691 : 1;
	24692 : 1;
	24693 : 1;
	24694 : 1;
	24695 : 1;
	24696 : 1;
	24697 : 1;
	24698 : 1;
	24699 : 1;
	24700 : 1;
	24701 : 1;
	24702 : 1;
	24703 : 1;
	24704 : 1;
	24705 : 1;
	24706 : 1;
	24707 : 1;
	24708 : 1;
	24709 : 1;
	24710 : 1;
	24711 : 1;
	24712 : 1;
	24713 : 1;
	24714 : 1;
	24715 : 1;
	24716 : 1;
	24717 : 1;
	24718 : 1;
	24719 : 1;
	24720 : 1;
	24721 : 1;
	24722 : 1;
	24723 : 1;
	24724 : 1;
	24725 : 1;
	24726 : 1;
	24727 : 1;
	24728 : 1;
	24729 : 1;
	24730 : 1;
	24731 : 1;
	24732 : 1;
	24733 : 1;
	24734 : 1;
	24735 : 1;
	24736 : 1;
	24737 : 1;
	24738 : 1;
	24739 : 1;
	24740 : 1;
	24741 : 1;
	24742 : 1;
	24743 : 1;
	24744 : 1;
	24745 : 1;
	24746 : 1;
	24747 : 1;
	24748 : 1;
	24749 : 1;
	24750 : 1;
	24751 : 1;
	24752 : 1;
	24753 : 1;
	24754 : 1;
	24755 : 1;
	24756 : 1;
	24757 : 1;
	24758 : 1;
	24759 : 1;
	24760 : 1;
	24761 : 1;
	24762 : 1;
	24763 : 1;
	24764 : 1;
	24765 : 1;
	24766 : 1;
	24767 : 1;
	24768 : 1;
	24769 : 1;
	24770 : 1;
	24771 : 1;
	24772 : 1;
	24773 : 1;
	24774 : 1;
	24775 : 1;
	24776 : 1;
	24777 : 1;
	24778 : 1;
	24779 : 1;
	24780 : 1;
	24781 : 1;
	24782 : 1;
	24783 : 1;
	24784 : 1;
	24785 : 1;
	24786 : 1;
	24787 : 1;
	24788 : 1;
	24789 : 1;
	24790 : 1;
	24791 : 1;
	24792 : 1;
	24793 : 1;
	24794 : 1;
	24795 : 1;
	24796 : 1;
	24797 : 1;
	24798 : 1;
	24799 : 1;
	24800 : 1;
	24801 : 1;
	24802 : 1;
	24803 : 1;
	24804 : 1;
	24805 : 1;
	24806 : 1;
	24807 : 1;
	24808 : 1;
	24809 : 1;
	24810 : 1;
	24811 : 1;
	24812 : 1;
	24813 : 1;
	24814 : 1;
	24815 : 1;
	24816 : 1;
	24817 : 1;
	24818 : 1;
	24819 : 1;
	24820 : 1;
	24821 : 1;
	24822 : 1;
	24823 : 1;
	24824 : 1;
	24825 : 1;
	24826 : 1;
	24827 : 1;
	24828 : 1;
	24829 : 1;
	24830 : 1;
	24831 : 1;
	24832 : 1;
	24833 : 1;
	24834 : 1;
	24835 : 1;
	24836 : 1;
	24837 : 1;
	24838 : 1;
	24839 : 1;
	24840 : 1;
	24841 : 1;
	24842 : 1;
	24843 : 1;
	24844 : 1;
	24845 : 1;
	24846 : 1;
	24847 : 1;
	24848 : 1;
	24849 : 1;
	24850 : 1;
	24851 : 1;
	24852 : 1;
	24853 : 1;
	24854 : 1;
	24855 : 1;
	24856 : 1;
	24857 : 1;
	24858 : 1;
	24859 : 1;
	24860 : 1;
	24861 : 1;
	24862 : 1;
	24863 : 1;
	24864 : 1;
	24865 : 1;
	24866 : 1;
	24867 : 1;
	24868 : 1;
	24869 : 1;
	24870 : 1;
	24871 : 1;
	24872 : 1;
	24873 : 1;
	24874 : 1;
	24875 : 1;
	24876 : 1;
	24877 : 1;
	24878 : 1;
	24879 : 1;
	24880 : 1;
	24881 : 1;
	24882 : 1;
	24883 : 1;
	24884 : 1;
	24885 : 1;
	24886 : 1;
	24887 : 1;
	24888 : 1;
	24889 : 1;
	24890 : 1;
	24891 : 1;
	24892 : 1;
	24893 : 1;
	24894 : 1;
	24895 : 1;
	24896 : 1;
	24897 : 1;
	24898 : 1;
	24899 : 1;
	24900 : 1;
	24901 : 1;
	24902 : 1;
	24903 : 1;
	24904 : 1;
	24905 : 1;
	24906 : 1;
	24907 : 1;
	24908 : 1;
	24909 : 1;
	24910 : 1;
	24911 : 1;
	24912 : 1;
	24913 : 1;
	24914 : 1;
	24915 : 1;
	24916 : 1;
	24917 : 1;
	24918 : 1;
	24919 : 1;
	24920 : 1;
	24921 : 1;
	24922 : 1;
	24923 : 1;
	24924 : 1;
	24925 : 1;
	24926 : 1;
	24927 : 1;
	24928 : 1;
	24929 : 1;
	24930 : 1;
	24931 : 1;
	24932 : 1;
	24933 : 1;
	24934 : 1;
	24935 : 1;
	24936 : 1;
	24937 : 1;
	24938 : 1;
	24939 : 1;
	24940 : 1;
	24941 : 1;
	24942 : 1;
	24943 : 1;
	24944 : 1;
	24945 : 1;
	24946 : 1;
	24947 : 1;
	24948 : 1;
	24949 : 1;
	24950 : 1;
	24951 : 1;
	24952 : 1;
	24953 : 1;
	24954 : 1;
	24955 : 1;
	24956 : 1;
	24957 : 1;
	24958 : 1;
	24959 : 1;
	24960 : 1;
	24961 : 1;
	24962 : 1;
	24963 : 1;
	24964 : 1;
	24965 : 1;
	24966 : 1;
	24967 : 1;
	24968 : 1;
	24969 : 1;
	24970 : 1;
	24971 : 1;
	24972 : 1;
	24973 : 1;
	24974 : 1;
	24975 : 1;
	24976 : 1;
	24977 : 1;
	24978 : 1;
	24979 : 1;
	24980 : 1;
	24981 : 1;
	24982 : 1;
	24983 : 1;
	24984 : 1;
	24985 : 1;
	24986 : 1;
	24987 : 1;
	24988 : 1;
	24989 : 1;
	24990 : 1;
	24991 : 1;
	24992 : 1;
	24993 : 1;
	24994 : 1;
	24995 : 1;
	24996 : 1;
	24997 : 1;
	24998 : 1;
	24999 : 1;
	25000 : 1;
	25001 : 1;
	25002 : 1;
	25003 : 1;
	25004 : 1;
	25005 : 1;
	25006 : 1;
	25007 : 1;
	25008 : 1;
	25009 : 1;
	25010 : 1;
	25011 : 1;
	25012 : 1;
	25013 : 1;
	25014 : 1;
	25015 : 1;
	25016 : 1;
	25017 : 1;
	25018 : 1;
	25019 : 1;
	25020 : 1;
	25021 : 1;
	25022 : 1;
	25023 : 1;
	25024 : 1;
	25025 : 1;
	25026 : 1;
	25027 : 1;
	25028 : 1;
	25029 : 1;
	25030 : 1;
	25031 : 1;
	25032 : 1;
	25033 : 1;
	25034 : 1;
	25035 : 1;
	25036 : 1;
	25037 : 1;
	25038 : 1;
	25039 : 1;
	25040 : 1;
	25041 : 1;
	25042 : 1;
	25043 : 1;
	25044 : 1;
	25045 : 1;
	25046 : 1;
	25047 : 1;
	25048 : 1;
	25049 : 1;
	25050 : 1;
	25051 : 1;
	25052 : 1;
	25053 : 1;
	25054 : 1;
	25055 : 1;
	25056 : 1;
	25057 : 1;
	25058 : 1;
	25059 : 1;
	25060 : 1;
	25061 : 1;
	25062 : 1;
	25063 : 1;
	25064 : 1;
	25065 : 1;
	25066 : 1;
	25067 : 1;
	25068 : 1;
	25069 : 1;
	25070 : 1;
	25071 : 1;
	25072 : 1;
	25073 : 1;
	25074 : 1;
	25075 : 1;
	25076 : 1;
	25077 : 1;
	25078 : 1;
	25079 : 1;
	25080 : 1;
	25081 : 1;
	25082 : 1;
	25083 : 1;
	25084 : 1;
	25085 : 1;
	25086 : 1;
	25087 : 1;
	25088 : 1;
	25089 : 1;
	25090 : 1;
	25091 : 1;
	25092 : 1;
	25093 : 1;
	25094 : 1;
	25095 : 1;
	25096 : 1;
	25097 : 1;
	25098 : 1;
	25099 : 1;
	25100 : 1;
	25101 : 1;
	25102 : 1;
	25103 : 1;
	25104 : 1;
	25105 : 1;
	25106 : 1;
	25107 : 1;
	25108 : 1;
	25109 : 1;
	25110 : 1;
	25111 : 1;
	25112 : 1;
	25113 : 1;
	25114 : 1;
	25115 : 1;
	25116 : 1;
	25117 : 1;
	25118 : 1;
	25119 : 1;
	25120 : 1;
	25121 : 1;
	25122 : 1;
	25123 : 1;
	25124 : 1;
	25125 : 1;
	25126 : 1;
	25127 : 1;
	25128 : 1;
	25129 : 1;
	25130 : 1;
	25131 : 1;
	25132 : 1;
	25133 : 1;
	25134 : 1;
	25135 : 1;
	25136 : 1;
	25137 : 1;
	25138 : 1;
	25139 : 1;
	25140 : 1;
	25141 : 1;
	25142 : 1;
	25143 : 1;
	25144 : 1;
	25145 : 1;
	25146 : 1;
	25147 : 1;
	25148 : 1;
	25149 : 1;
	25150 : 1;
	25151 : 1;
	25152 : 1;
	25153 : 1;
	25154 : 1;
	25155 : 1;
	25156 : 1;
	25157 : 1;
	25158 : 1;
	25159 : 1;
	25160 : 1;
	25161 : 1;
	25162 : 1;
	25163 : 1;
	25164 : 1;
	25165 : 1;
	25166 : 1;
	25167 : 1;
	25168 : 1;
	25169 : 1;
	25170 : 1;
	25171 : 1;
	25172 : 1;
	25173 : 1;
	25174 : 1;
	25175 : 1;
	25176 : 1;
	25177 : 1;
	25178 : 1;
	25179 : 1;
	25180 : 1;
	25181 : 1;
	25182 : 1;
	25183 : 1;
	25184 : 1;
	25185 : 1;
	25186 : 1;
	25187 : 1;
	25188 : 1;
	25189 : 1;
	25190 : 1;
	25191 : 1;
	25192 : 1;
	25193 : 1;
	25194 : 1;
	25195 : 1;
	25196 : 1;
	25197 : 1;
	25198 : 1;
	25199 : 1;
	25200 : 1;
	25201 : 1;
	25202 : 1;
	25203 : 1;
	25204 : 1;
	25205 : 1;
	25206 : 1;
	25207 : 1;
	25208 : 1;
	25209 : 1;
	25210 : 1;
	25211 : 1;
	25212 : 1;
	25213 : 1;
	25214 : 1;
	25215 : 1;
	25216 : 1;
	25217 : 1;
	25218 : 1;
	25219 : 1;
	25220 : 1;
	25221 : 1;
	25222 : 1;
	25223 : 1;
	25224 : 1;
	25225 : 1;
	25226 : 1;
	25227 : 1;
	25228 : 1;
	25229 : 1;
	25230 : 1;
	25231 : 1;
	25232 : 1;
	25233 : 1;
	25234 : 1;
	25235 : 1;
	25236 : 1;
	25237 : 1;
	25238 : 1;
	25239 : 1;
	25240 : 1;
	25241 : 1;
	25242 : 1;
	25243 : 1;
	25244 : 1;
	25245 : 1;
	25246 : 1;
	25247 : 1;
	25248 : 1;
	25249 : 1;
	25250 : 1;
	25251 : 1;
	25252 : 1;
	25253 : 1;
	25254 : 1;
	25255 : 1;
	25256 : 1;
	25257 : 1;
	25258 : 1;
	25259 : 1;
	25260 : 1;
	25261 : 1;
	25262 : 1;
	25263 : 1;
	25264 : 1;
	25265 : 1;
	25266 : 1;
	25267 : 1;
	25268 : 1;
	25269 : 1;
	25270 : 1;
	25271 : 1;
	25272 : 1;
	25273 : 1;
	25274 : 1;
	25275 : 1;
	25276 : 1;
	25277 : 1;
	25278 : 1;
	25279 : 1;
	25280 : 1;
	25281 : 1;
	25282 : 1;
	25283 : 1;
	25284 : 1;
	25285 : 1;
	25286 : 1;
	25287 : 1;
	25288 : 1;
	25289 : 1;
	25290 : 1;
	25291 : 1;
	25292 : 1;
	25293 : 1;
	25294 : 1;
	25295 : 0;
	25296 : 0;
	25297 : 1;
	25298 : 1;
	25299 : 1;
	25300 : 1;
	25301 : 1;
	25302 : 1;
	25303 : 1;
	25304 : 1;
	25305 : 1;
	25306 : 1;
	25307 : 1;
	25308 : 1;
	25309 : 1;
	25310 : 1;
	25311 : 1;
	25312 : 1;
	25313 : 1;
	25314 : 1;
	25315 : 1;
	25316 : 1;
	25317 : 1;
	25318 : 1;
	25319 : 1;
	25320 : 1;
	25321 : 1;
	25322 : 1;
	25323 : 1;
	25324 : 1;
	25325 : 1;
	25326 : 1;
	25327 : 1;
	25328 : 1;
	25329 : 1;
	25330 : 1;
	25331 : 1;
	25332 : 1;
	25333 : 1;
	25334 : 1;
	25335 : 1;
	25336 : 1;
	25337 : 1;
	25338 : 1;
	25339 : 1;
	25340 : 1;
	25341 : 1;
	25342 : 1;
	25343 : 1;
	25344 : 1;
	25345 : 1;
	25346 : 1;
	25347 : 1;
	25348 : 1;
	25349 : 1;
	25350 : 1;
	25351 : 1;
	25352 : 1;
	25353 : 1;
	25354 : 1;
	25355 : 1;
	25356 : 1;
	25357 : 1;
	25358 : 1;
	25359 : 1;
	25360 : 1;
	25361 : 1;
	25362 : 1;
	25363 : 1;
	25364 : 1;
	25365 : 1;
	25366 : 1;
	25367 : 1;
	25368 : 1;
	25369 : 1;
	25370 : 1;
	25371 : 1;
	25372 : 1;
	25373 : 1;
	25374 : 1;
	25375 : 1;
	25376 : 1;
	25377 : 1;
	25378 : 1;
	25379 : 1;
	25380 : 1;
	25381 : 1;
	25382 : 1;
	25383 : 1;
	25384 : 1;
	25385 : 1;
	25386 : 1;
	25387 : 1;
	25388 : 1;
	25389 : 1;
	25390 : 1;
	25391 : 1;
	25392 : 1;
	25393 : 1;
	25394 : 1;
	25395 : 1;
	25396 : 1;
	25397 : 1;
	25398 : 1;
	25399 : 1;
	25400 : 1;
	25401 : 1;
	25402 : 1;
	25403 : 1;
	25404 : 1;
	25405 : 1;
	25406 : 1;
	25407 : 1;
	25408 : 1;
	25409 : 1;
	25410 : 1;
	25411 : 1;
	25412 : 1;
	25413 : 1;
	25414 : 1;
	25415 : 1;
	25416 : 1;
	25417 : 1;
	25418 : 1;
	25419 : 1;
	25420 : 1;
	25421 : 1;
	25422 : 1;
	25423 : 1;
	25424 : 1;
	25425 : 1;
	25426 : 1;
	25427 : 1;
	25428 : 1;
	25429 : 1;
	25430 : 1;
	25431 : 1;
	25432 : 1;
	25433 : 1;
	25434 : 1;
	25435 : 1;
	25436 : 1;
	25437 : 1;
	25438 : 1;
	25439 : 1;
	25440 : 1;
	25441 : 1;
	25442 : 1;
	25443 : 1;
	25444 : 1;
	25445 : 1;
	25446 : 1;
	25447 : 1;
	25448 : 1;
	25449 : 1;
	25450 : 1;
	25451 : 1;
	25452 : 1;
	25453 : 1;
	25454 : 1;
	25455 : 1;
	25456 : 1;
	25457 : 1;
	25458 : 1;
	25459 : 1;
	25460 : 1;
	25461 : 1;
	25462 : 1;
	25463 : 1;
	25464 : 1;
	25465 : 1;
	25466 : 1;
	25467 : 1;
	25468 : 1;
	25469 : 1;
	25470 : 1;
	25471 : 1;
	25472 : 1;
	25473 : 1;
	25474 : 1;
	25475 : 1;
	25476 : 1;
	25477 : 1;
	25478 : 1;
	25479 : 1;
	25480 : 1;
	25481 : 1;
	25482 : 1;
	25483 : 1;
	25484 : 1;
	25485 : 1;
	25486 : 1;
	25487 : 1;
	25488 : 1;
	25489 : 1;
	25490 : 1;
	25491 : 1;
	25492 : 1;
	25493 : 1;
	25494 : 1;
	25495 : 1;
	25496 : 1;
	25497 : 1;
	25498 : 1;
	25499 : 1;
	25500 : 1;
	25501 : 1;
	25502 : 1;
	25503 : 1;
	25504 : 1;
	25505 : 1;
	25506 : 1;
	25507 : 1;
	25508 : 1;
	25509 : 1;
	25510 : 1;
	25511 : 1;
	25512 : 1;
	25513 : 1;
	25514 : 1;
	25515 : 1;
	25516 : 1;
	25517 : 1;
	25518 : 1;
	25519 : 1;
	25520 : 1;
	25521 : 1;
	25522 : 1;
	25523 : 1;
	25524 : 1;
	25525 : 1;
	25526 : 1;
	25527 : 1;
	25528 : 1;
	25529 : 1;
	25530 : 1;
	25531 : 1;
	25532 : 1;
	25533 : 1;
	25534 : 1;
	25535 : 0;
	25536 : 0;
	25537 : 1;
	25538 : 1;
	25539 : 1;
	25540 : 1;
	25541 : 1;
	25542 : 1;
	25543 : 1;
	25544 : 1;
	25545 : 1;
	25546 : 1;
	25547 : 1;
	25548 : 1;
	25549 : 1;
	25550 : 1;
	25551 : 1;
	25552 : 1;
	25553 : 1;
	25554 : 1;
	25555 : 1;
	25556 : 1;
	25557 : 1;
	25558 : 1;
	25559 : 1;
	25560 : 1;
	25561 : 1;
	25562 : 1;
	25563 : 1;
	25564 : 1;
	25565 : 1;
	25566 : 1;
	25567 : 1;
	25568 : 1;
	25569 : 1;
	25570 : 1;
	25571 : 1;
	25572 : 1;
	25573 : 1;
	25574 : 1;
	25575 : 1;
	25576 : 1;
	25577 : 1;
	25578 : 1;
	25579 : 1;
	25580 : 1;
	25581 : 1;
	25582 : 1;
	25583 : 1;
	25584 : 1;
	25585 : 1;
	25586 : 1;
	25587 : 1;
	25588 : 1;
	25589 : 1;
	25590 : 1;
	25591 : 1;
	25592 : 1;
	25593 : 1;
	25594 : 1;
	25595 : 1;
	25596 : 1;
	25597 : 1;
	25598 : 1;
	25599 : 1;
	25600 : 1;
	25601 : 1;
	25602 : 1;
	25603 : 1;
	25604 : 1;
	25605 : 1;
	25606 : 1;
	25607 : 1;
	25608 : 1;
	25609 : 1;
	25610 : 1;
	25611 : 1;
	25612 : 1;
	25613 : 1;
	25614 : 1;
	25615 : 1;
	25616 : 1;
	25617 : 1;
	25618 : 1;
	25619 : 1;
	25620 : 1;
	25621 : 1;
	25622 : 1;
	25623 : 1;
	25624 : 1;
	25625 : 1;
	25626 : 1;
	25627 : 1;
	25628 : 1;
	25629 : 1;
	25630 : 1;
	25631 : 1;
	25632 : 1;
	25633 : 1;
	25634 : 1;
	25635 : 1;
	25636 : 1;
	25637 : 1;
	25638 : 1;
	25639 : 1;
	25640 : 1;
	25641 : 1;
	25642 : 1;
	25643 : 1;
	25644 : 1;
	25645 : 1;
	25646 : 1;
	25647 : 1;
	25648 : 1;
	25649 : 1;
	25650 : 1;
	25651 : 1;
	25652 : 1;
	25653 : 1;
	25654 : 1;
	25655 : 1;
	25656 : 1;
	25657 : 1;
	25658 : 1;
	25659 : 1;
	25660 : 1;
	25661 : 1;
	25662 : 1;
	25663 : 1;
	25664 : 1;
	25665 : 1;
	25666 : 1;
	25667 : 1;
	25668 : 1;
	25669 : 1;
	25670 : 1;
	25671 : 1;
	25672 : 1;
	25673 : 1;
	25674 : 1;
	25675 : 1;
	25676 : 1;
	25677 : 1;
	25678 : 1;
	25679 : 1;
	25680 : 1;
	25681 : 1;
	25682 : 1;
	25683 : 1;
	25684 : 1;
	25685 : 1;
	25686 : 1;
	25687 : 1;
	25688 : 1;
	25689 : 1;
	25690 : 1;
	25691 : 1;
	25692 : 1;
	25693 : 1;
	25694 : 1;
	25695 : 1;
	25696 : 1;
	25697 : 1;
	25698 : 1;
	25699 : 1;
	25700 : 1;
	25701 : 1;
	25702 : 1;
	25703 : 1;
	25704 : 1;
	25705 : 1;
	25706 : 1;
	25707 : 1;
	25708 : 1;
	25709 : 1;
	25710 : 1;
	25711 : 1;
	25712 : 1;
	25713 : 1;
	25714 : 1;
	25715 : 1;
	25716 : 1;
	25717 : 1;
	25718 : 1;
	25719 : 1;
	25720 : 1;
	25721 : 1;
	25722 : 1;
	25723 : 1;
	25724 : 1;
	25725 : 1;
	25726 : 1;
	25727 : 1;
	25728 : 1;
	25729 : 1;
	25730 : 1;
	25731 : 1;
	25732 : 1;
	25733 : 1;
	25734 : 1;
	25735 : 1;
	25736 : 1;
	25737 : 1;
	25738 : 1;
	25739 : 1;
	25740 : 1;
	25741 : 1;
	25742 : 1;
	25743 : 1;
	25744 : 1;
	25745 : 1;
	25746 : 1;
	25747 : 1;
	25748 : 1;
	25749 : 1;
	25750 : 1;
	25751 : 1;
	25752 : 1;
	25753 : 1;
	25754 : 1;
	25755 : 1;
	25756 : 1;
	25757 : 1;
	25758 : 1;
	25759 : 1;
	25760 : 1;
	25761 : 1;
	25762 : 1;
	25763 : 1;
	25764 : 1;
	25765 : 1;
	25766 : 1;
	25767 : 1;
	25768 : 1;
	25769 : 1;
	25770 : 1;
	25771 : 1;
	25772 : 1;
	25773 : 1;
	25774 : 1;
	25775 : 0;
	25776 : 0;
	25777 : 1;
	25778 : 1;
	25779 : 1;
	25780 : 1;
	25781 : 1;
	25782 : 1;
	25783 : 1;
	25784 : 1;
	25785 : 1;
	25786 : 1;
	25787 : 1;
	25788 : 1;
	25789 : 1;
	25790 : 1;
	25791 : 1;
	25792 : 1;
	25793 : 1;
	25794 : 1;
	25795 : 1;
	25796 : 1;
	25797 : 1;
	25798 : 1;
	25799 : 1;
	25800 : 1;
	25801 : 1;
	25802 : 1;
	25803 : 1;
	25804 : 1;
	25805 : 1;
	25806 : 1;
	25807 : 1;
	25808 : 1;
	25809 : 1;
	25810 : 1;
	25811 : 1;
	25812 : 1;
	25813 : 1;
	25814 : 1;
	25815 : 1;
	25816 : 1;
	25817 : 1;
	25818 : 1;
	25819 : 1;
	25820 : 1;
	25821 : 1;
	25822 : 1;
	25823 : 1;
	25824 : 1;
	25825 : 1;
	25826 : 1;
	25827 : 1;
	25828 : 1;
	25829 : 1;
	25830 : 1;
	25831 : 1;
	25832 : 1;
	25833 : 1;
	25834 : 1;
	25835 : 1;
	25836 : 1;
	25837 : 1;
	25838 : 1;
	25839 : 1;
	25840 : 1;
	25841 : 1;
	25842 : 1;
	25843 : 1;
	25844 : 1;
	25845 : 1;
	25846 : 1;
	25847 : 1;
	25848 : 1;
	25849 : 1;
	25850 : 1;
	25851 : 1;
	25852 : 1;
	25853 : 1;
	25854 : 1;
	25855 : 1;
	25856 : 1;
	25857 : 1;
	25858 : 1;
	25859 : 1;
	25860 : 1;
	25861 : 1;
	25862 : 1;
	25863 : 1;
	25864 : 1;
	25865 : 1;
	25866 : 1;
	25867 : 1;
	25868 : 1;
	25869 : 1;
	25870 : 1;
	25871 : 1;
	25872 : 1;
	25873 : 1;
	25874 : 1;
	25875 : 1;
	25876 : 1;
	25877 : 1;
	25878 : 1;
	25879 : 1;
	25880 : 1;
	25881 : 1;
	25882 : 1;
	25883 : 1;
	25884 : 1;
	25885 : 1;
	25886 : 1;
	25887 : 1;
	25888 : 1;
	25889 : 1;
	25890 : 1;
	25891 : 1;
	25892 : 1;
	25893 : 1;
	25894 : 1;
	25895 : 1;
	25896 : 1;
	25897 : 1;
	25898 : 1;
	25899 : 1;
	25900 : 1;
	25901 : 1;
	25902 : 1;
	25903 : 1;
	25904 : 1;
	25905 : 1;
	25906 : 1;
	25907 : 1;
	25908 : 1;
	25909 : 1;
	25910 : 1;
	25911 : 1;
	25912 : 1;
	25913 : 1;
	25914 : 1;
	25915 : 1;
	25916 : 1;
	25917 : 1;
	25918 : 1;
	25919 : 1;
	25920 : 1;
	25921 : 1;
	25922 : 1;
	25923 : 1;
	25924 : 1;
	25925 : 1;
	25926 : 1;
	25927 : 1;
	25928 : 1;
	25929 : 1;
	25930 : 1;
	25931 : 1;
	25932 : 1;
	25933 : 1;
	25934 : 1;
	25935 : 1;
	25936 : 1;
	25937 : 1;
	25938 : 1;
	25939 : 1;
	25940 : 1;
	25941 : 1;
	25942 : 1;
	25943 : 1;
	25944 : 1;
	25945 : 1;
	25946 : 1;
	25947 : 1;
	25948 : 1;
	25949 : 1;
	25950 : 1;
	25951 : 1;
	25952 : 1;
	25953 : 1;
	25954 : 1;
	25955 : 1;
	25956 : 1;
	25957 : 1;
	25958 : 1;
	25959 : 1;
	25960 : 1;
	25961 : 1;
	25962 : 1;
	25963 : 1;
	25964 : 1;
	25965 : 1;
	25966 : 1;
	25967 : 1;
	25968 : 1;
	25969 : 1;
	25970 : 1;
	25971 : 1;
	25972 : 1;
	25973 : 1;
	25974 : 1;
	25975 : 1;
	25976 : 1;
	25977 : 1;
	25978 : 1;
	25979 : 1;
	25980 : 1;
	25981 : 1;
	25982 : 1;
	25983 : 1;
	25984 : 1;
	25985 : 1;
	25986 : 1;
	25987 : 1;
	25988 : 1;
	25989 : 1;
	25990 : 1;
	25991 : 1;
	25992 : 1;
	25993 : 1;
	25994 : 1;
	25995 : 1;
	25996 : 1;
	25997 : 1;
	25998 : 1;
	25999 : 1;
	26000 : 1;
	26001 : 1;
	26002 : 1;
	26003 : 1;
	26004 : 1;
	26005 : 1;
	26006 : 1;
	26007 : 1;
	26008 : 1;
	26009 : 1;
	26010 : 1;
	26011 : 1;
	26012 : 1;
	26013 : 1;
	26014 : 1;
	26015 : 0;
	26016 : 0;
	26017 : 1;
	26018 : 1;
	26019 : 1;
	26020 : 1;
	26021 : 1;
	26022 : 1;
	26023 : 1;
	26024 : 1;
	26025 : 1;
	26026 : 1;
	26027 : 1;
	26028 : 1;
	26029 : 1;
	26030 : 1;
	26031 : 1;
	26032 : 1;
	26033 : 1;
	26034 : 1;
	26035 : 1;
	26036 : 1;
	26037 : 1;
	26038 : 1;
	26039 : 1;
	26040 : 1;
	26041 : 1;
	26042 : 1;
	26043 : 1;
	26044 : 1;
	26045 : 1;
	26046 : 1;
	26047 : 1;
	26048 : 1;
	26049 : 1;
	26050 : 1;
	26051 : 1;
	26052 : 1;
	26053 : 1;
	26054 : 1;
	26055 : 1;
	26056 : 1;
	26057 : 1;
	26058 : 1;
	26059 : 1;
	26060 : 1;
	26061 : 1;
	26062 : 1;
	26063 : 1;
	26064 : 1;
	26065 : 1;
	26066 : 1;
	26067 : 1;
	26068 : 1;
	26069 : 1;
	26070 : 1;
	26071 : 1;
	26072 : 1;
	26073 : 1;
	26074 : 1;
	26075 : 1;
	26076 : 1;
	26077 : 1;
	26078 : 1;
	26079 : 1;
	26080 : 1;
	26081 : 1;
	26082 : 1;
	26083 : 1;
	26084 : 1;
	26085 : 1;
	26086 : 1;
	26087 : 1;
	26088 : 1;
	26089 : 1;
	26090 : 1;
	26091 : 1;
	26092 : 1;
	26093 : 1;
	26094 : 1;
	26095 : 1;
	26096 : 1;
	26097 : 1;
	26098 : 1;
	26099 : 1;
	26100 : 1;
	26101 : 1;
	26102 : 1;
	26103 : 1;
	26104 : 1;
	26105 : 1;
	26106 : 1;
	26107 : 1;
	26108 : 1;
	26109 : 1;
	26110 : 1;
	26111 : 1;
	26112 : 1;
	26113 : 1;
	26114 : 1;
	26115 : 1;
	26116 : 1;
	26117 : 1;
	26118 : 1;
	26119 : 1;
	26120 : 1;
	26121 : 1;
	26122 : 1;
	26123 : 1;
	26124 : 1;
	26125 : 1;
	26126 : 1;
	26127 : 1;
	26128 : 1;
	26129 : 1;
	26130 : 1;
	26131 : 1;
	26132 : 1;
	26133 : 1;
	26134 : 1;
	26135 : 1;
	26136 : 1;
	26137 : 1;
	26138 : 1;
	26139 : 1;
	26140 : 1;
	26141 : 1;
	26142 : 1;
	26143 : 1;
	26144 : 1;
	26145 : 1;
	26146 : 1;
	26147 : 1;
	26148 : 1;
	26149 : 1;
	26150 : 1;
	26151 : 1;
	26152 : 1;
	26153 : 1;
	26154 : 1;
	26155 : 1;
	26156 : 1;
	26157 : 1;
	26158 : 1;
	26159 : 1;
	26160 : 1;
	26161 : 1;
	26162 : 1;
	26163 : 1;
	26164 : 1;
	26165 : 1;
	26166 : 1;
	26167 : 1;
	26168 : 1;
	26169 : 1;
	26170 : 1;
	26171 : 1;
	26172 : 1;
	26173 : 1;
	26174 : 1;
	26175 : 1;
	26176 : 1;
	26177 : 1;
	26178 : 1;
	26179 : 1;
	26180 : 1;
	26181 : 1;
	26182 : 1;
	26183 : 1;
	26184 : 1;
	26185 : 1;
	26186 : 1;
	26187 : 1;
	26188 : 1;
	26189 : 1;
	26190 : 1;
	26191 : 1;
	26192 : 1;
	26193 : 1;
	26194 : 1;
	26195 : 1;
	26196 : 1;
	26197 : 1;
	26198 : 1;
	26199 : 1;
	26200 : 1;
	26201 : 1;
	26202 : 1;
	26203 : 1;
	26204 : 1;
	26205 : 1;
	26206 : 1;
	26207 : 1;
	26208 : 1;
	26209 : 1;
	26210 : 1;
	26211 : 1;
	26212 : 1;
	26213 : 1;
	26214 : 1;
	26215 : 1;
	26216 : 1;
	26217 : 1;
	26218 : 1;
	26219 : 1;
	26220 : 1;
	26221 : 1;
	26222 : 1;
	26223 : 1;
	26224 : 1;
	26225 : 1;
	26226 : 1;
	26227 : 1;
	26228 : 1;
	26229 : 1;
	26230 : 1;
	26231 : 1;
	26232 : 1;
	26233 : 1;
	26234 : 1;
	26235 : 1;
	26236 : 1;
	26237 : 1;
	26238 : 1;
	26239 : 1;
	26240 : 1;
	26241 : 1;
	26242 : 1;
	26243 : 1;
	26244 : 1;
	26245 : 1;
	26246 : 1;
	26247 : 1;
	26248 : 1;
	26249 : 1;
	26250 : 1;
	26251 : 1;
	26252 : 1;
	26253 : 1;
	26254 : 1;
	26255 : 0;
	26256 : 1;
	26257 : 1;
	26258 : 1;
	26259 : 1;
	26260 : 1;
	26261 : 1;
	26262 : 1;
	26263 : 1;
	26264 : 1;
	26265 : 1;
	26266 : 1;
	26267 : 1;
	26268 : 1;
	26269 : 1;
	26270 : 1;
	26271 : 1;
	26272 : 1;
	26273 : 1;
	26274 : 1;
	26275 : 1;
	26276 : 1;
	26277 : 1;
	26278 : 1;
	26279 : 1;
	26280 : 1;
	26281 : 1;
	26282 : 1;
	26283 : 1;
	26284 : 1;
	26285 : 1;
	26286 : 1;
	26287 : 1;
	26288 : 1;
	26289 : 1;
	26290 : 1;
	26291 : 1;
	26292 : 1;
	26293 : 1;
	26294 : 1;
	26295 : 1;
	26296 : 1;
	26297 : 1;
	26298 : 1;
	26299 : 1;
	26300 : 1;
	26301 : 1;
	26302 : 1;
	26303 : 1;
	26304 : 1;
	26305 : 1;
	26306 : 1;
	26307 : 1;
	26308 : 1;
	26309 : 1;
	26310 : 1;
	26311 : 1;
	26312 : 1;
	26313 : 1;
	26314 : 1;
	26315 : 1;
	26316 : 1;
	26317 : 1;
	26318 : 1;
	26319 : 1;
	26320 : 1;
	26321 : 1;
	26322 : 1;
	26323 : 1;
	26324 : 1;
	26325 : 1;
	26326 : 1;
	26327 : 1;
	26328 : 1;
	26329 : 1;
	26330 : 1;
	26331 : 1;
	26332 : 1;
	26333 : 1;
	26334 : 1;
	26335 : 1;
	26336 : 1;
	26337 : 1;
	26338 : 1;
	26339 : 1;
	26340 : 1;
	26341 : 1;
	26342 : 1;
	26343 : 1;
	26344 : 1;
	26345 : 1;
	26346 : 1;
	26347 : 1;
	26348 : 1;
	26349 : 1;
	26350 : 1;
	26351 : 1;
	26352 : 1;
	26353 : 1;
	26354 : 1;
	26355 : 1;
	26356 : 1;
	26357 : 1;
	26358 : 1;
	26359 : 1;
	26360 : 1;
	26361 : 1;
	26362 : 1;
	26363 : 1;
	26364 : 1;
	26365 : 1;
	26366 : 1;
	26367 : 1;
	26368 : 1;
	26369 : 1;
	26370 : 1;
	26371 : 1;
	26372 : 1;
	26373 : 1;
	26374 : 1;
	26375 : 1;
	26376 : 1;
	26377 : 1;
	26378 : 1;
	26379 : 1;
	26380 : 1;
	26381 : 1;
	26382 : 1;
	26383 : 1;
	26384 : 1;
	26385 : 1;
	26386 : 1;
	26387 : 1;
	26388 : 1;
	26389 : 1;
	26390 : 1;
	26391 : 1;
	26392 : 1;
	26393 : 1;
	26394 : 1;
	26395 : 1;
	26396 : 1;
	26397 : 1;
	26398 : 1;
	26399 : 1;
	26400 : 1;
	26401 : 1;
	26402 : 1;
	26403 : 1;
	26404 : 1;
	26405 : 1;
	26406 : 1;
	26407 : 1;
	26408 : 1;
	26409 : 1;
	26410 : 1;
	26411 : 1;
	26412 : 1;
	26413 : 1;
	26414 : 1;
	26415 : 1;
	26416 : 1;
	26417 : 1;
	26418 : 1;
	26419 : 1;
	26420 : 0;
	26421 : 0;
	26422 : 0;
	26423 : 0;
	26424 : 1;
	26425 : 1;
	26426 : 1;
	26427 : 1;
	26428 : 1;
	26429 : 1;
	26430 : 1;
	26431 : 1;
	26432 : 1;
	26433 : 1;
	26434 : 1;
	26435 : 1;
	26436 : 1;
	26437 : 1;
	26438 : 1;
	26439 : 1;
	26440 : 1;
	26441 : 1;
	26442 : 1;
	26443 : 1;
	26444 : 1;
	26445 : 1;
	26446 : 1;
	26447 : 1;
	26448 : 1;
	26449 : 1;
	26450 : 1;
	26451 : 1;
	26452 : 1;
	26453 : 1;
	26454 : 1;
	26455 : 1;
	26456 : 1;
	26457 : 1;
	26458 : 1;
	26459 : 1;
	26460 : 1;
	26461 : 1;
	26462 : 1;
	26463 : 1;
	26464 : 1;
	26465 : 1;
	26466 : 1;
	26467 : 0;
	26468 : 1;
	26469 : 1;
	26470 : 1;
	26471 : 0;
	26472 : 0;
	26473 : 1;
	26474 : 1;
	26475 : 1;
	26476 : 1;
	26477 : 1;
	26478 : 1;
	26479 : 1;
	26480 : 1;
	26481 : 1;
	26482 : 1;
	26483 : 1;
	26484 : 1;
	26485 : 1;
	26486 : 1;
	26487 : 1;
	26488 : 1;
	26489 : 1;
	26490 : 1;
	26491 : 1;
	26492 : 1;
	26493 : 1;
	26494 : 1;
	26495 : 1;
	26496 : 1;
	26497 : 1;
	26498 : 1;
	26499 : 1;
	26500 : 1;
	26501 : 1;
	26502 : 1;
	26503 : 1;
	26504 : 1;
	26505 : 1;
	26506 : 1;
	26507 : 1;
	26508 : 1;
	26509 : 1;
	26510 : 1;
	26511 : 1;
	26512 : 1;
	26513 : 1;
	26514 : 1;
	26515 : 1;
	26516 : 1;
	26517 : 1;
	26518 : 1;
	26519 : 1;
	26520 : 1;
	26521 : 1;
	26522 : 1;
	26523 : 1;
	26524 : 1;
	26525 : 1;
	26526 : 1;
	26527 : 1;
	26528 : 1;
	26529 : 1;
	26530 : 1;
	26531 : 1;
	26532 : 1;
	26533 : 1;
	26534 : 0;
	26535 : 1;
	26536 : 1;
	26537 : 1;
	26538 : 1;
	26539 : 1;
	26540 : 1;
	26541 : 1;
	26542 : 1;
	26543 : 1;
	26544 : 1;
	26545 : 1;
	26546 : 1;
	26547 : 1;
	26548 : 1;
	26549 : 1;
	26550 : 1;
	26551 : 1;
	26552 : 1;
	26553 : 1;
	26554 : 1;
	26555 : 1;
	26556 : 1;
	26557 : 1;
	26558 : 1;
	26559 : 1;
	26560 : 1;
	26561 : 1;
	26562 : 1;
	26563 : 1;
	26564 : 1;
	26565 : 1;
	26566 : 1;
	26567 : 1;
	26568 : 1;
	26569 : 1;
	26570 : 1;
	26571 : 1;
	26572 : 1;
	26573 : 1;
	26574 : 1;
	26575 : 1;
	26576 : 1;
	26577 : 1;
	26578 : 1;
	26579 : 1;
	26580 : 1;
	26581 : 1;
	26582 : 1;
	26583 : 1;
	26584 : 1;
	26585 : 1;
	26586 : 1;
	26587 : 1;
	26588 : 1;
	26589 : 1;
	26590 : 0;
	26591 : 1;
	26592 : 1;
	26593 : 1;
	26594 : 0;
	26595 : 1;
	26596 : 1;
	26597 : 1;
	26598 : 1;
	26599 : 1;
	26600 : 1;
	26601 : 1;
	26602 : 1;
	26603 : 1;
	26604 : 1;
	26605 : 1;
	26606 : 1;
	26607 : 1;
	26608 : 1;
	26609 : 1;
	26610 : 1;
	26611 : 1;
	26612 : 1;
	26613 : 1;
	26614 : 1;
	26615 : 1;
	26616 : 1;
	26617 : 1;
	26618 : 1;
	26619 : 1;
	26620 : 1;
	26621 : 1;
	26622 : 1;
	26623 : 1;
	26624 : 1;
	26625 : 1;
	26626 : 1;
	26627 : 1;
	26628 : 1;
	26629 : 1;
	26630 : 1;
	26631 : 1;
	26632 : 1;
	26633 : 1;
	26634 : 1;
	26635 : 1;
	26636 : 1;
	26637 : 1;
	26638 : 1;
	26639 : 1;
	26640 : 1;
	26641 : 1;
	26642 : 1;
	26643 : 1;
	26644 : 1;
	26645 : 1;
	26646 : 1;
	26647 : 1;
	26648 : 1;
	26649 : 1;
	26650 : 1;
	26651 : 1;
	26652 : 1;
	26653 : 1;
	26654 : 1;
	26655 : 1;
	26656 : 1;
	26657 : 1;
	26658 : 1;
	26659 : 0;
	26660 : 1;
	26661 : 1;
	26662 : 1;
	26663 : 0;
	26664 : 1;
	26665 : 1;
	26666 : 1;
	26667 : 1;
	26668 : 1;
	26669 : 1;
	26670 : 1;
	26671 : 1;
	26672 : 1;
	26673 : 1;
	26674 : 1;
	26675 : 1;
	26676 : 1;
	26677 : 1;
	26678 : 1;
	26679 : 1;
	26680 : 1;
	26681 : 1;
	26682 : 1;
	26683 : 1;
	26684 : 1;
	26685 : 1;
	26686 : 1;
	26687 : 1;
	26688 : 1;
	26689 : 1;
	26690 : 1;
	26691 : 1;
	26692 : 1;
	26693 : 1;
	26694 : 1;
	26695 : 0;
	26696 : 0;
	26697 : 1;
	26698 : 1;
	26699 : 1;
	26700 : 1;
	26701 : 1;
	26702 : 1;
	26703 : 1;
	26704 : 1;
	26705 : 1;
	26706 : 1;
	26707 : 1;
	26708 : 1;
	26709 : 1;
	26710 : 0;
	26711 : 1;
	26712 : 1;
	26713 : 1;
	26714 : 1;
	26715 : 1;
	26716 : 1;
	26717 : 1;
	26718 : 1;
	26719 : 1;
	26720 : 1;
	26721 : 1;
	26722 : 1;
	26723 : 1;
	26724 : 1;
	26725 : 1;
	26726 : 1;
	26727 : 1;
	26728 : 1;
	26729 : 1;
	26730 : 1;
	26731 : 1;
	26732 : 1;
	26733 : 1;
	26734 : 1;
	26735 : 1;
	26736 : 1;
	26737 : 1;
	26738 : 1;
	26739 : 1;
	26740 : 1;
	26741 : 1;
	26742 : 1;
	26743 : 1;
	26744 : 1;
	26745 : 1;
	26746 : 1;
	26747 : 1;
	26748 : 1;
	26749 : 1;
	26750 : 1;
	26751 : 1;
	26752 : 1;
	26753 : 1;
	26754 : 1;
	26755 : 1;
	26756 : 1;
	26757 : 1;
	26758 : 1;
	26759 : 1;
	26760 : 1;
	26761 : 1;
	26762 : 1;
	26763 : 1;
	26764 : 1;
	26765 : 1;
	26766 : 1;
	26767 : 1;
	26768 : 1;
	26769 : 1;
	26770 : 1;
	26771 : 1;
	26772 : 1;
	26773 : 1;
	26774 : 0;
	26775 : 1;
	26776 : 1;
	26777 : 1;
	26778 : 1;
	26779 : 1;
	26780 : 1;
	26781 : 1;
	26782 : 1;
	26783 : 1;
	26784 : 1;
	26785 : 1;
	26786 : 1;
	26787 : 1;
	26788 : 1;
	26789 : 0;
	26790 : 1;
	26791 : 1;
	26792 : 1;
	26793 : 1;
	26794 : 1;
	26795 : 1;
	26796 : 1;
	26797 : 1;
	26798 : 1;
	26799 : 1;
	26800 : 1;
	26801 : 1;
	26802 : 1;
	26803 : 1;
	26804 : 1;
	26805 : 1;
	26806 : 1;
	26807 : 1;
	26808 : 1;
	26809 : 1;
	26810 : 1;
	26811 : 1;
	26812 : 1;
	26813 : 1;
	26814 : 1;
	26815 : 1;
	26816 : 1;
	26817 : 1;
	26818 : 1;
	26819 : 1;
	26820 : 1;
	26821 : 1;
	26822 : 1;
	26823 : 1;
	26824 : 1;
	26825 : 1;
	26826 : 1;
	26827 : 1;
	26828 : 1;
	26829 : 1;
	26830 : 0;
	26831 : 1;
	26832 : 1;
	26833 : 1;
	26834 : 0;
	26835 : 1;
	26836 : 1;
	26837 : 1;
	26838 : 1;
	26839 : 1;
	26840 : 1;
	26841 : 1;
	26842 : 1;
	26843 : 1;
	26844 : 1;
	26845 : 1;
	26846 : 1;
	26847 : 1;
	26848 : 1;
	26849 : 1;
	26850 : 1;
	26851 : 1;
	26852 : 1;
	26853 : 1;
	26854 : 1;
	26855 : 1;
	26856 : 1;
	26857 : 1;
	26858 : 1;
	26859 : 1;
	26860 : 1;
	26861 : 1;
	26862 : 1;
	26863 : 1;
	26864 : 1;
	26865 : 1;
	26866 : 1;
	26867 : 1;
	26868 : 1;
	26869 : 1;
	26870 : 1;
	26871 : 1;
	26872 : 1;
	26873 : 1;
	26874 : 1;
	26875 : 1;
	26876 : 1;
	26877 : 1;
	26878 : 1;
	26879 : 1;
	26880 : 1;
	26881 : 1;
	26882 : 1;
	26883 : 1;
	26884 : 1;
	26885 : 1;
	26886 : 1;
	26887 : 1;
	26888 : 1;
	26889 : 1;
	26890 : 1;
	26891 : 1;
	26892 : 1;
	26893 : 1;
	26894 : 1;
	26895 : 1;
	26896 : 1;
	26897 : 1;
	26898 : 1;
	26899 : 0;
	26900 : 1;
	26901 : 1;
	26902 : 1;
	26903 : 1;
	26904 : 1;
	26905 : 1;
	26906 : 1;
	26907 : 1;
	26908 : 1;
	26909 : 1;
	26910 : 1;
	26911 : 1;
	26912 : 1;
	26913 : 1;
	26914 : 1;
	26915 : 1;
	26916 : 1;
	26917 : 1;
	26918 : 1;
	26919 : 1;
	26920 : 1;
	26921 : 1;
	26922 : 1;
	26923 : 1;
	26924 : 1;
	26925 : 1;
	26926 : 1;
	26927 : 1;
	26928 : 1;
	26929 : 1;
	26930 : 1;
	26931 : 1;
	26932 : 1;
	26933 : 1;
	26934 : 1;
	26935 : 0;
	26936 : 0;
	26937 : 1;
	26938 : 1;
	26939 : 1;
	26940 : 1;
	26941 : 1;
	26942 : 1;
	26943 : 1;
	26944 : 1;
	26945 : 1;
	26946 : 1;
	26947 : 1;
	26948 : 1;
	26949 : 1;
	26950 : 0;
	26951 : 1;
	26952 : 1;
	26953 : 1;
	26954 : 1;
	26955 : 1;
	26956 : 1;
	26957 : 1;
	26958 : 1;
	26959 : 1;
	26960 : 1;
	26961 : 1;
	26962 : 1;
	26963 : 1;
	26964 : 1;
	26965 : 1;
	26966 : 1;
	26967 : 1;
	26968 : 1;
	26969 : 1;
	26970 : 1;
	26971 : 1;
	26972 : 1;
	26973 : 1;
	26974 : 1;
	26975 : 1;
	26976 : 1;
	26977 : 1;
	26978 : 1;
	26979 : 1;
	26980 : 1;
	26981 : 1;
	26982 : 1;
	26983 : 1;
	26984 : 1;
	26985 : 1;
	26986 : 1;
	26987 : 1;
	26988 : 1;
	26989 : 1;
	26990 : 1;
	26991 : 1;
	26992 : 1;
	26993 : 1;
	26994 : 1;
	26995 : 1;
	26996 : 1;
	26997 : 1;
	26998 : 1;
	26999 : 1;
	27000 : 1;
	27001 : 1;
	27002 : 1;
	27003 : 1;
	27004 : 1;
	27005 : 1;
	27006 : 1;
	27007 : 1;
	27008 : 1;
	27009 : 1;
	27010 : 1;
	27011 : 1;
	27012 : 1;
	27013 : 0;
	27014 : 0;
	27015 : 1;
	27016 : 1;
	27017 : 1;
	27018 : 1;
	27019 : 1;
	27020 : 1;
	27021 : 1;
	27022 : 1;
	27023 : 1;
	27024 : 1;
	27025 : 1;
	27026 : 1;
	27027 : 1;
	27028 : 1;
	27029 : 0;
	27030 : 0;
	27031 : 1;
	27032 : 1;
	27033 : 1;
	27034 : 1;
	27035 : 1;
	27036 : 1;
	27037 : 1;
	27038 : 1;
	27039 : 1;
	27040 : 1;
	27041 : 1;
	27042 : 1;
	27043 : 1;
	27044 : 1;
	27045 : 1;
	27046 : 1;
	27047 : 1;
	27048 : 1;
	27049 : 1;
	27050 : 1;
	27051 : 1;
	27052 : 1;
	27053 : 1;
	27054 : 1;
	27055 : 1;
	27056 : 1;
	27057 : 1;
	27058 : 1;
	27059 : 1;
	27060 : 1;
	27061 : 1;
	27062 : 1;
	27063 : 1;
	27064 : 1;
	27065 : 1;
	27066 : 1;
	27067 : 1;
	27068 : 1;
	27069 : 1;
	27070 : 0;
	27071 : 1;
	27072 : 1;
	27073 : 1;
	27074 : 0;
	27075 : 1;
	27076 : 1;
	27077 : 1;
	27078 : 1;
	27079 : 1;
	27080 : 1;
	27081 : 1;
	27082 : 1;
	27083 : 1;
	27084 : 1;
	27085 : 1;
	27086 : 1;
	27087 : 1;
	27088 : 1;
	27089 : 1;
	27090 : 1;
	27091 : 1;
	27092 : 1;
	27093 : 1;
	27094 : 1;
	27095 : 1;
	27096 : 1;
	27097 : 1;
	27098 : 1;
	27099 : 1;
	27100 : 1;
	27101 : 1;
	27102 : 1;
	27103 : 1;
	27104 : 1;
	27105 : 1;
	27106 : 1;
	27107 : 1;
	27108 : 1;
	27109 : 1;
	27110 : 1;
	27111 : 1;
	27112 : 1;
	27113 : 1;
	27114 : 1;
	27115 : 1;
	27116 : 1;
	27117 : 1;
	27118 : 1;
	27119 : 1;
	27120 : 1;
	27121 : 1;
	27122 : 1;
	27123 : 1;
	27124 : 1;
	27125 : 1;
	27126 : 1;
	27127 : 1;
	27128 : 1;
	27129 : 1;
	27130 : 1;
	27131 : 1;
	27132 : 1;
	27133 : 1;
	27134 : 1;
	27135 : 1;
	27136 : 1;
	27137 : 1;
	27138 : 1;
	27139 : 0;
	27140 : 1;
	27141 : 1;
	27142 : 1;
	27143 : 1;
	27144 : 1;
	27145 : 1;
	27146 : 0;
	27147 : 0;
	27148 : 0;
	27149 : 0;
	27150 : 1;
	27151 : 0;
	27152 : 0;
	27153 : 0;
	27154 : 0;
	27155 : 1;
	27156 : 1;
	27157 : 0;
	27158 : 0;
	27159 : 0;
	27160 : 0;
	27161 : 1;
	27162 : 1;
	27163 : 0;
	27164 : 1;
	27165 : 0;
	27166 : 0;
	27167 : 1;
	27168 : 1;
	27169 : 0;
	27170 : 0;
	27171 : 0;
	27172 : 0;
	27173 : 0;
	27174 : 1;
	27175 : 0;
	27176 : 0;
	27177 : 0;
	27178 : 0;
	27179 : 1;
	27180 : 0;
	27181 : 0;
	27182 : 0;
	27183 : 0;
	27184 : 1;
	27185 : 1;
	27186 : 1;
	27187 : 0;
	27188 : 1;
	27189 : 0;
	27190 : 0;
	27191 : 0;
	27192 : 0;
	27193 : 1;
	27194 : 1;
	27195 : 1;
	27196 : 0;
	27197 : 1;
	27198 : 1;
	27199 : 1;
	27200 : 0;
	27201 : 0;
	27202 : 1;
	27203 : 0;
	27204 : 0;
	27205 : 0;
	27206 : 0;
	27207 : 1;
	27208 : 1;
	27209 : 0;
	27210 : 1;
	27211 : 1;
	27212 : 0;
	27213 : 1;
	27214 : 1;
	27215 : 1;
	27216 : 1;
	27217 : 1;
	27218 : 0;
	27219 : 0;
	27220 : 0;
	27221 : 0;
	27222 : 1;
	27223 : 1;
	27224 : 0;
	27225 : 0;
	27226 : 0;
	27227 : 0;
	27228 : 1;
	27229 : 1;
	27230 : 1;
	27231 : 1;
	27232 : 0;
	27233 : 0;
	27234 : 0;
	27235 : 0;
	27236 : 1;
	27237 : 1;
	27238 : 0;
	27239 : 1;
	27240 : 0;
	27241 : 0;
	27242 : 1;
	27243 : 1;
	27244 : 0;
	27245 : 0;
	27246 : 0;
	27247 : 0;
	27248 : 0;
	27249 : 1;
	27250 : 0;
	27251 : 0;
	27252 : 0;
	27253 : 0;
	27254 : 0;
	27255 : 1;
	27256 : 0;
	27257 : 1;
	27258 : 1;
	27259 : 0;
	27260 : 1;
	27261 : 1;
	27262 : 1;
	27263 : 0;
	27264 : 0;
	27265 : 0;
	27266 : 0;
	27267 : 1;
	27268 : 0;
	27269 : 0;
	27270 : 0;
	27271 : 0;
	27272 : 1;
	27273 : 0;
	27274 : 0;
	27275 : 0;
	27276 : 0;
	27277 : 0;
	27278 : 0;
	27279 : 1;
	27280 : 1;
	27281 : 0;
	27282 : 0;
	27283 : 0;
	27284 : 0;
	27285 : 1;
	27286 : 1;
	27287 : 1;
	27288 : 1;
	27289 : 1;
	27290 : 1;
	27291 : 1;
	27292 : 1;
	27293 : 1;
	27294 : 1;
	27295 : 0;
	27296 : 0;
	27297 : 0;
	27298 : 0;
	27299 : 0;
	27300 : 0;
	27301 : 0;
	27302 : 0;
	27303 : 0;
	27304 : 1;
	27305 : 1;
	27306 : 0;
	27307 : 0;
	27308 : 0;
	27309 : 0;
	27310 : 0;
	27311 : 1;
	27312 : 1;
	27313 : 1;
	27314 : 0;
	27315 : 0;
	27316 : 0;
	27317 : 0;
	27318 : 0;
	27319 : 1;
	27320 : 1;
	27321 : 0;
	27322 : 0;
	27323 : 0;
	27324 : 0;
	27325 : 0;
	27326 : 0;
	27327 : 0;
	27328 : 1;
	27329 : 1;
	27330 : 1;
	27331 : 0;
	27332 : 1;
	27333 : 0;
	27334 : 0;
	27335 : 0;
	27336 : 0;
	27337 : 1;
	27338 : 1;
	27339 : 1;
	27340 : 1;
	27341 : 1;
	27342 : 1;
	27343 : 1;
	27344 : 1;
	27345 : 1;
	27346 : 1;
	27347 : 1;
	27348 : 1;
	27349 : 1;
	27350 : 1;
	27351 : 1;
	27352 : 1;
	27353 : 1;
	27354 : 1;
	27355 : 1;
	27356 : 1;
	27357 : 1;
	27358 : 1;
	27359 : 1;
	27360 : 1;
	27361 : 1;
	27362 : 1;
	27363 : 1;
	27364 : 1;
	27365 : 1;
	27366 : 1;
	27367 : 1;
	27368 : 1;
	27369 : 1;
	27370 : 1;
	27371 : 1;
	27372 : 1;
	27373 : 1;
	27374 : 1;
	27375 : 1;
	27376 : 1;
	27377 : 1;
	27378 : 1;
	27379 : 0;
	27380 : 1;
	27381 : 1;
	27382 : 1;
	27383 : 1;
	27384 : 1;
	27385 : 0;
	27386 : 1;
	27387 : 1;
	27388 : 1;
	27389 : 0;
	27390 : 0;
	27391 : 0;
	27392 : 0;
	27393 : 1;
	27394 : 0;
	27395 : 0;
	27396 : 1;
	27397 : 0;
	27398 : 1;
	27399 : 1;
	27400 : 1;
	27401 : 0;
	27402 : 1;
	27403 : 0;
	27404 : 0;
	27405 : 1;
	27406 : 1;
	27407 : 1;
	27408 : 0;
	27409 : 1;
	27410 : 1;
	27411 : 1;
	27412 : 0;
	27413 : 0;
	27414 : 1;
	27415 : 0;
	27416 : 0;
	27417 : 1;
	27418 : 1;
	27419 : 1;
	27420 : 0;
	27421 : 1;
	27422 : 1;
	27423 : 1;
	27424 : 1;
	27425 : 1;
	27426 : 1;
	27427 : 0;
	27428 : 1;
	27429 : 1;
	27430 : 0;
	27431 : 1;
	27432 : 1;
	27433 : 1;
	27434 : 1;
	27435 : 1;
	27436 : 0;
	27437 : 1;
	27438 : 1;
	27439 : 1;
	27440 : 0;
	27441 : 0;
	27442 : 0;
	27443 : 0;
	27444 : 1;
	27445 : 1;
	27446 : 1;
	27447 : 0;
	27448 : 1;
	27449 : 0;
	27450 : 1;
	27451 : 1;
	27452 : 0;
	27453 : 1;
	27454 : 1;
	27455 : 1;
	27456 : 1;
	27457 : 1;
	27458 : 0;
	27459 : 0;
	27460 : 1;
	27461 : 1;
	27462 : 1;
	27463 : 0;
	27464 : 0;
	27465 : 1;
	27466 : 1;
	27467 : 0;
	27468 : 0;
	27469 : 1;
	27470 : 1;
	27471 : 1;
	27472 : 0;
	27473 : 1;
	27474 : 1;
	27475 : 1;
	27476 : 0;
	27477 : 1;
	27478 : 0;
	27479 : 0;
	27480 : 1;
	27481 : 1;
	27482 : 1;
	27483 : 0;
	27484 : 1;
	27485 : 1;
	27486 : 1;
	27487 : 0;
	27488 : 0;
	27489 : 0;
	27490 : 0;
	27491 : 1;
	27492 : 1;
	27493 : 1;
	27494 : 0;
	27495 : 1;
	27496 : 0;
	27497 : 1;
	27498 : 1;
	27499 : 0;
	27500 : 1;
	27501 : 1;
	27502 : 0;
	27503 : 1;
	27504 : 1;
	27505 : 1;
	27506 : 0;
	27507 : 1;
	27508 : 1;
	27509 : 0;
	27510 : 1;
	27511 : 1;
	27512 : 1;
	27513 : 0;
	27514 : 0;
	27515 : 0;
	27516 : 0;
	27517 : 1;
	27518 : 0;
	27519 : 0;
	27520 : 1;
	27521 : 0;
	27522 : 1;
	27523 : 1;
	27524 : 1;
	27525 : 0;
	27526 : 1;
	27527 : 1;
	27528 : 1;
	27529 : 1;
	27530 : 1;
	27531 : 1;
	27532 : 1;
	27533 : 1;
	27534 : 0;
	27535 : 1;
	27536 : 1;
	27537 : 1;
	27538 : 0;
	27539 : 0;
	27540 : 0;
	27541 : 0;
	27542 : 1;
	27543 : 0;
	27544 : 0;
	27545 : 1;
	27546 : 0;
	27547 : 1;
	27548 : 1;
	27549 : 1;
	27550 : 0;
	27551 : 1;
	27552 : 1;
	27553 : 1;
	27554 : 0;
	27555 : 1;
	27556 : 1;
	27557 : 1;
	27558 : 0;
	27559 : 1;
	27560 : 0;
	27561 : 1;
	27562 : 1;
	27563 : 1;
	27564 : 0;
	27565 : 0;
	27566 : 0;
	27567 : 0;
	27568 : 1;
	27569 : 1;
	27570 : 0;
	27571 : 0;
	27572 : 1;
	27573 : 0;
	27574 : 1;
	27575 : 1;
	27576 : 1;
	27577 : 0;
	27578 : 1;
	27579 : 1;
	27580 : 1;
	27581 : 1;
	27582 : 1;
	27583 : 1;
	27584 : 1;
	27585 : 1;
	27586 : 1;
	27587 : 1;
	27588 : 1;
	27589 : 1;
	27590 : 1;
	27591 : 1;
	27592 : 1;
	27593 : 1;
	27594 : 1;
	27595 : 1;
	27596 : 1;
	27597 : 1;
	27598 : 1;
	27599 : 1;
	27600 : 1;
	27601 : 1;
	27602 : 1;
	27603 : 1;
	27604 : 1;
	27605 : 1;
	27606 : 1;
	27607 : 1;
	27608 : 1;
	27609 : 1;
	27610 : 1;
	27611 : 1;
	27612 : 1;
	27613 : 1;
	27614 : 1;
	27615 : 1;
	27616 : 1;
	27617 : 1;
	27618 : 1;
	27619 : 0;
	27620 : 1;
	27621 : 1;
	27622 : 1;
	27623 : 1;
	27624 : 1;
	27625 : 0;
	27626 : 1;
	27627 : 1;
	27628 : 1;
	27629 : 0;
	27630 : 0;
	27631 : 0;
	27632 : 0;
	27633 : 1;
	27634 : 0;
	27635 : 0;
	27636 : 1;
	27637 : 0;
	27638 : 1;
	27639 : 1;
	27640 : 1;
	27641 : 0;
	27642 : 1;
	27643 : 0;
	27644 : 1;
	27645 : 1;
	27646 : 1;
	27647 : 1;
	27648 : 0;
	27649 : 1;
	27650 : 1;
	27651 : 1;
	27652 : 0;
	27653 : 0;
	27654 : 1;
	27655 : 0;
	27656 : 0;
	27657 : 1;
	27658 : 1;
	27659 : 1;
	27660 : 1;
	27661 : 0;
	27662 : 0;
	27663 : 1;
	27664 : 1;
	27665 : 1;
	27666 : 1;
	27667 : 0;
	27668 : 1;
	27669 : 1;
	27670 : 0;
	27671 : 1;
	27672 : 1;
	27673 : 1;
	27674 : 1;
	27675 : 1;
	27676 : 0;
	27677 : 1;
	27678 : 1;
	27679 : 1;
	27680 : 0;
	27681 : 0;
	27682 : 0;
	27683 : 0;
	27684 : 1;
	27685 : 1;
	27686 : 1;
	27687 : 0;
	27688 : 1;
	27689 : 0;
	27690 : 1;
	27691 : 1;
	27692 : 0;
	27693 : 1;
	27694 : 1;
	27695 : 1;
	27696 : 1;
	27697 : 1;
	27698 : 0;
	27699 : 1;
	27700 : 1;
	27701 : 1;
	27702 : 1;
	27703 : 0;
	27704 : 0;
	27705 : 0;
	27706 : 0;
	27707 : 0;
	27708 : 0;
	27709 : 1;
	27710 : 1;
	27711 : 1;
	27712 : 0;
	27713 : 1;
	27714 : 1;
	27715 : 1;
	27716 : 0;
	27717 : 1;
	27718 : 0;
	27719 : 1;
	27720 : 1;
	27721 : 1;
	27722 : 1;
	27723 : 0;
	27724 : 1;
	27725 : 1;
	27726 : 1;
	27727 : 0;
	27728 : 0;
	27729 : 0;
	27730 : 0;
	27731 : 1;
	27732 : 1;
	27733 : 1;
	27734 : 0;
	27735 : 1;
	27736 : 0;
	27737 : 1;
	27738 : 1;
	27739 : 0;
	27740 : 1;
	27741 : 1;
	27742 : 0;
	27743 : 1;
	27744 : 1;
	27745 : 1;
	27746 : 0;
	27747 : 1;
	27748 : 1;
	27749 : 0;
	27750 : 1;
	27751 : 1;
	27752 : 1;
	27753 : 0;
	27754 : 0;
	27755 : 0;
	27756 : 0;
	27757 : 1;
	27758 : 0;
	27759 : 0;
	27760 : 1;
	27761 : 0;
	27762 : 1;
	27763 : 1;
	27764 : 1;
	27765 : 0;
	27766 : 1;
	27767 : 1;
	27768 : 1;
	27769 : 1;
	27770 : 1;
	27771 : 1;
	27772 : 1;
	27773 : 1;
	27774 : 0;
	27775 : 1;
	27776 : 1;
	27777 : 1;
	27778 : 0;
	27779 : 0;
	27780 : 0;
	27781 : 0;
	27782 : 1;
	27783 : 0;
	27784 : 0;
	27785 : 1;
	27786 : 0;
	27787 : 1;
	27788 : 1;
	27789 : 1;
	27790 : 0;
	27791 : 1;
	27792 : 1;
	27793 : 1;
	27794 : 0;
	27795 : 1;
	27796 : 1;
	27797 : 1;
	27798 : 0;
	27799 : 1;
	27800 : 0;
	27801 : 1;
	27802 : 1;
	27803 : 1;
	27804 : 0;
	27805 : 0;
	27806 : 1;
	27807 : 0;
	27808 : 0;
	27809 : 0;
	27810 : 0;
	27811 : 1;
	27812 : 1;
	27813 : 0;
	27814 : 0;
	27815 : 0;
	27816 : 0;
	27817 : 0;
	27818 : 1;
	27819 : 1;
	27820 : 1;
	27821 : 1;
	27822 : 1;
	27823 : 1;
	27824 : 1;
	27825 : 1;
	27826 : 1;
	27827 : 1;
	27828 : 1;
	27829 : 1;
	27830 : 1;
	27831 : 1;
	27832 : 1;
	27833 : 1;
	27834 : 1;
	27835 : 1;
	27836 : 1;
	27837 : 1;
	27838 : 1;
	27839 : 1;
	27840 : 1;
	27841 : 1;
	27842 : 1;
	27843 : 1;
	27844 : 1;
	27845 : 1;
	27846 : 1;
	27847 : 1;
	27848 : 1;
	27849 : 1;
	27850 : 1;
	27851 : 1;
	27852 : 1;
	27853 : 1;
	27854 : 1;
	27855 : 1;
	27856 : 1;
	27857 : 1;
	27858 : 1;
	27859 : 0;
	27860 : 1;
	27861 : 1;
	27862 : 1;
	27863 : 0;
	27864 : 1;
	27865 : 0;
	27866 : 1;
	27867 : 1;
	27868 : 1;
	27869 : 0;
	27870 : 0;
	27871 : 0;
	27872 : 0;
	27873 : 1;
	27874 : 0;
	27875 : 0;
	27876 : 1;
	27877 : 0;
	27878 : 1;
	27879 : 1;
	27880 : 1;
	27881 : 0;
	27882 : 1;
	27883 : 0;
	27884 : 1;
	27885 : 1;
	27886 : 1;
	27887 : 1;
	27888 : 0;
	27889 : 1;
	27890 : 1;
	27891 : 0;
	27892 : 0;
	27893 : 0;
	27894 : 1;
	27895 : 0;
	27896 : 0;
	27897 : 1;
	27898 : 1;
	27899 : 1;
	27900 : 1;
	27901 : 1;
	27902 : 1;
	27903 : 0;
	27904 : 1;
	27905 : 1;
	27906 : 1;
	27907 : 0;
	27908 : 1;
	27909 : 1;
	27910 : 0;
	27911 : 1;
	27912 : 1;
	27913 : 1;
	27914 : 1;
	27915 : 1;
	27916 : 0;
	27917 : 1;
	27918 : 1;
	27919 : 1;
	27920 : 0;
	27921 : 0;
	27922 : 0;
	27923 : 0;
	27924 : 1;
	27925 : 1;
	27926 : 1;
	27927 : 0;
	27928 : 1;
	27929 : 0;
	27930 : 1;
	27931 : 1;
	27932 : 0;
	27933 : 1;
	27934 : 1;
	27935 : 1;
	27936 : 1;
	27937 : 1;
	27938 : 0;
	27939 : 1;
	27940 : 1;
	27941 : 1;
	27942 : 1;
	27943 : 0;
	27944 : 0;
	27945 : 1;
	27946 : 1;
	27947 : 1;
	27948 : 1;
	27949 : 1;
	27950 : 1;
	27951 : 1;
	27952 : 0;
	27953 : 1;
	27954 : 1;
	27955 : 1;
	27956 : 0;
	27957 : 1;
	27958 : 0;
	27959 : 1;
	27960 : 1;
	27961 : 1;
	27962 : 1;
	27963 : 0;
	27964 : 1;
	27965 : 1;
	27966 : 0;
	27967 : 0;
	27968 : 0;
	27969 : 0;
	27970 : 0;
	27971 : 1;
	27972 : 1;
	27973 : 1;
	27974 : 0;
	27975 : 1;
	27976 : 0;
	27977 : 1;
	27978 : 1;
	27979 : 0;
	27980 : 1;
	27981 : 1;
	27982 : 0;
	27983 : 1;
	27984 : 1;
	27985 : 0;
	27986 : 0;
	27987 : 1;
	27988 : 1;
	27989 : 0;
	27990 : 1;
	27991 : 1;
	27992 : 1;
	27993 : 0;
	27994 : 0;
	27995 : 0;
	27996 : 0;
	27997 : 1;
	27998 : 0;
	27999 : 0;
	28000 : 1;
	28001 : 0;
	28002 : 1;
	28003 : 1;
	28004 : 1;
	28005 : 0;
	28006 : 1;
	28007 : 0;
	28008 : 0;
	28009 : 1;
	28010 : 1;
	28011 : 1;
	28012 : 1;
	28013 : 1;
	28014 : 0;
	28015 : 1;
	28016 : 1;
	28017 : 0;
	28018 : 0;
	28019 : 0;
	28020 : 0;
	28021 : 0;
	28022 : 1;
	28023 : 0;
	28024 : 0;
	28025 : 1;
	28026 : 0;
	28027 : 1;
	28028 : 1;
	28029 : 1;
	28030 : 0;
	28031 : 1;
	28032 : 1;
	28033 : 1;
	28034 : 0;
	28035 : 1;
	28036 : 1;
	28037 : 1;
	28038 : 0;
	28039 : 1;
	28040 : 0;
	28041 : 1;
	28042 : 1;
	28043 : 0;
	28044 : 0;
	28045 : 0;
	28046 : 1;
	28047 : 0;
	28048 : 0;
	28049 : 0;
	28050 : 0;
	28051 : 1;
	28052 : 1;
	28053 : 0;
	28054 : 1;
	28055 : 1;
	28056 : 1;
	28057 : 1;
	28058 : 1;
	28059 : 1;
	28060 : 1;
	28061 : 1;
	28062 : 1;
	28063 : 1;
	28064 : 1;
	28065 : 1;
	28066 : 1;
	28067 : 1;
	28068 : 1;
	28069 : 1;
	28070 : 1;
	28071 : 1;
	28072 : 1;
	28073 : 1;
	28074 : 1;
	28075 : 1;
	28076 : 1;
	28077 : 1;
	28078 : 1;
	28079 : 1;
	28080 : 1;
	28081 : 1;
	28082 : 1;
	28083 : 1;
	28084 : 1;
	28085 : 1;
	28086 : 1;
	28087 : 1;
	28088 : 1;
	28089 : 1;
	28090 : 1;
	28091 : 1;
	28092 : 1;
	28093 : 1;
	28094 : 1;
	28095 : 1;
	28096 : 1;
	28097 : 1;
	28098 : 1;
	28099 : 1;
	28100 : 0;
	28101 : 0;
	28102 : 0;
	28103 : 1;
	28104 : 1;
	28105 : 1;
	28106 : 0;
	28107 : 0;
	28108 : 0;
	28109 : 0;
	28110 : 1;
	28111 : 0;
	28112 : 0;
	28113 : 1;
	28114 : 0;
	28115 : 0;
	28116 : 1;
	28117 : 1;
	28118 : 0;
	28119 : 0;
	28120 : 0;
	28121 : 0;
	28122 : 1;
	28123 : 0;
	28124 : 1;
	28125 : 1;
	28126 : 1;
	28127 : 1;
	28128 : 1;
	28129 : 0;
	28130 : 0;
	28131 : 0;
	28132 : 0;
	28133 : 0;
	28134 : 1;
	28135 : 0;
	28136 : 0;
	28137 : 0;
	28138 : 0;
	28139 : 1;
	28140 : 0;
	28141 : 0;
	28142 : 0;
	28143 : 0;
	28144 : 1;
	28145 : 1;
	28146 : 1;
	28147 : 0;
	28148 : 1;
	28149 : 1;
	28150 : 0;
	28151 : 1;
	28152 : 1;
	28153 : 1;
	28154 : 1;
	28155 : 1;
	28156 : 1;
	28157 : 0;
	28158 : 0;
	28159 : 0;
	28160 : 0;
	28161 : 0;
	28162 : 1;
	28163 : 0;
	28164 : 0;
	28165 : 0;
	28166 : 0;
	28167 : 1;
	28168 : 1;
	28169 : 1;
	28170 : 0;
	28171 : 0;
	28172 : 1;
	28173 : 0;
	28174 : 1;
	28175 : 1;
	28176 : 1;
	28177 : 1;
	28178 : 0;
	28179 : 1;
	28180 : 1;
	28181 : 1;
	28182 : 1;
	28183 : 1;
	28184 : 0;
	28185 : 0;
	28186 : 0;
	28187 : 0;
	28188 : 0;
	28189 : 1;
	28190 : 1;
	28191 : 1;
	28192 : 1;
	28193 : 0;
	28194 : 0;
	28195 : 0;
	28196 : 0;
	28197 : 1;
	28198 : 0;
	28199 : 1;
	28200 : 1;
	28201 : 1;
	28202 : 1;
	28203 : 1;
	28204 : 0;
	28205 : 0;
	28206 : 0;
	28207 : 0;
	28208 : 0;
	28209 : 1;
	28210 : 0;
	28211 : 0;
	28212 : 0;
	28213 : 0;
	28214 : 0;
	28215 : 1;
	28216 : 1;
	28217 : 0;
	28218 : 0;
	28219 : 1;
	28220 : 0;
	28221 : 1;
	28222 : 1;
	28223 : 0;
	28224 : 0;
	28225 : 1;
	28226 : 0;
	28227 : 1;
	28228 : 1;
	28229 : 0;
	28230 : 0;
	28231 : 0;
	28232 : 0;
	28233 : 0;
	28234 : 0;
	28235 : 0;
	28236 : 0;
	28237 : 1;
	28238 : 0;
	28239 : 0;
	28240 : 1;
	28241 : 1;
	28242 : 0;
	28243 : 0;
	28244 : 0;
	28245 : 0;
	28246 : 1;
	28247 : 0;
	28248 : 0;
	28249 : 1;
	28250 : 1;
	28251 : 1;
	28252 : 1;
	28253 : 1;
	28254 : 1;
	28255 : 0;
	28256 : 0;
	28257 : 0;
	28258 : 0;
	28259 : 0;
	28260 : 0;
	28261 : 0;
	28262 : 1;
	28263 : 0;
	28264 : 0;
	28265 : 1;
	28266 : 1;
	28267 : 0;
	28268 : 0;
	28269 : 0;
	28270 : 0;
	28271 : 1;
	28272 : 1;
	28273 : 1;
	28274 : 0;
	28275 : 1;
	28276 : 1;
	28277 : 1;
	28278 : 0;
	28279 : 1;
	28280 : 1;
	28281 : 0;
	28282 : 0;
	28283 : 0;
	28284 : 0;
	28285 : 0;
	28286 : 1;
	28287 : 1;
	28288 : 0;
	28289 : 0;
	28290 : 1;
	28291 : 1;
	28292 : 1;
	28293 : 1;
	28294 : 0;
	28295 : 0;
	28296 : 0;
	28297 : 0;
	28298 : 1;
	28299 : 1;
	28300 : 1;
	28301 : 1;
	28302 : 1;
	28303 : 1;
	28304 : 1;
	28305 : 1;
	28306 : 1;
	28307 : 1;
	28308 : 1;
	28309 : 1;
	28310 : 1;
	28311 : 1;
	28312 : 1;
	28313 : 1;
	28314 : 1;
	28315 : 1;
	28316 : 1;
	28317 : 1;
	28318 : 1;
	28319 : 1;
	28320 : 1;
	28321 : 1;
	28322 : 1;
	28323 : 1;
	28324 : 1;
	28325 : 1;
	28326 : 1;
	28327 : 1;
	28328 : 1;
	28329 : 1;
	28330 : 1;
	28331 : 1;
	28332 : 1;
	28333 : 1;
	28334 : 1;
	28335 : 1;
	28336 : 1;
	28337 : 1;
	28338 : 1;
	28339 : 1;
	28340 : 1;
	28341 : 1;
	28342 : 1;
	28343 : 1;
	28344 : 1;
	28345 : 1;
	28346 : 1;
	28347 : 1;
	28348 : 1;
	28349 : 1;
	28350 : 1;
	28351 : 1;
	28352 : 1;
	28353 : 1;
	28354 : 1;
	28355 : 1;
	28356 : 1;
	28357 : 1;
	28358 : 1;
	28359 : 1;
	28360 : 1;
	28361 : 0;
	28362 : 1;
	28363 : 1;
	28364 : 1;
	28365 : 1;
	28366 : 1;
	28367 : 1;
	28368 : 1;
	28369 : 1;
	28370 : 1;
	28371 : 1;
	28372 : 1;
	28373 : 1;
	28374 : 1;
	28375 : 1;
	28376 : 1;
	28377 : 1;
	28378 : 1;
	28379 : 1;
	28380 : 1;
	28381 : 1;
	28382 : 1;
	28383 : 1;
	28384 : 1;
	28385 : 1;
	28386 : 1;
	28387 : 1;
	28388 : 1;
	28389 : 1;
	28390 : 1;
	28391 : 1;
	28392 : 1;
	28393 : 1;
	28394 : 1;
	28395 : 1;
	28396 : 1;
	28397 : 1;
	28398 : 1;
	28399 : 1;
	28400 : 0;
	28401 : 0;
	28402 : 1;
	28403 : 1;
	28404 : 1;
	28405 : 1;
	28406 : 1;
	28407 : 1;
	28408 : 1;
	28409 : 1;
	28410 : 1;
	28411 : 1;
	28412 : 1;
	28413 : 1;
	28414 : 1;
	28415 : 1;
	28416 : 1;
	28417 : 1;
	28418 : 1;
	28419 : 1;
	28420 : 1;
	28421 : 1;
	28422 : 1;
	28423 : 1;
	28424 : 1;
	28425 : 1;
	28426 : 1;
	28427 : 1;
	28428 : 1;
	28429 : 1;
	28430 : 1;
	28431 : 1;
	28432 : 1;
	28433 : 1;
	28434 : 1;
	28435 : 1;
	28436 : 0;
	28437 : 1;
	28438 : 1;
	28439 : 1;
	28440 : 1;
	28441 : 1;
	28442 : 1;
	28443 : 1;
	28444 : 1;
	28445 : 1;
	28446 : 1;
	28447 : 1;
	28448 : 1;
	28449 : 1;
	28450 : 1;
	28451 : 1;
	28452 : 1;
	28453 : 1;
	28454 : 1;
	28455 : 1;
	28456 : 1;
	28457 : 1;
	28458 : 1;
	28459 : 1;
	28460 : 1;
	28461 : 1;
	28462 : 1;
	28463 : 1;
	28464 : 1;
	28465 : 1;
	28466 : 1;
	28467 : 1;
	28468 : 1;
	28469 : 1;
	28470 : 1;
	28471 : 1;
	28472 : 1;
	28473 : 1;
	28474 : 1;
	28475 : 1;
	28476 : 1;
	28477 : 1;
	28478 : 1;
	28479 : 1;
	28480 : 1;
	28481 : 1;
	28482 : 1;
	28483 : 1;
	28484 : 1;
	28485 : 0;
	28486 : 1;
	28487 : 1;
	28488 : 0;
	28489 : 1;
	28490 : 1;
	28491 : 1;
	28492 : 1;
	28493 : 1;
	28494 : 1;
	28495 : 1;
	28496 : 1;
	28497 : 1;
	28498 : 1;
	28499 : 1;
	28500 : 1;
	28501 : 1;
	28502 : 1;
	28503 : 1;
	28504 : 1;
	28505 : 1;
	28506 : 1;
	28507 : 1;
	28508 : 1;
	28509 : 1;
	28510 : 1;
	28511 : 1;
	28512 : 1;
	28513 : 1;
	28514 : 1;
	28515 : 1;
	28516 : 1;
	28517 : 1;
	28518 : 1;
	28519 : 1;
	28520 : 1;
	28521 : 1;
	28522 : 1;
	28523 : 1;
	28524 : 1;
	28525 : 1;
	28526 : 1;
	28527 : 1;
	28528 : 1;
	28529 : 1;
	28530 : 1;
	28531 : 1;
	28532 : 1;
	28533 : 1;
	28534 : 1;
	28535 : 1;
	28536 : 1;
	28537 : 1;
	28538 : 1;
	28539 : 1;
	28540 : 1;
	28541 : 1;
	28542 : 1;
	28543 : 1;
	28544 : 1;
	28545 : 1;
	28546 : 1;
	28547 : 1;
	28548 : 1;
	28549 : 1;
	28550 : 1;
	28551 : 1;
	28552 : 1;
	28553 : 1;
	28554 : 1;
	28555 : 1;
	28556 : 1;
	28557 : 1;
	28558 : 1;
	28559 : 1;
	28560 : 1;
	28561 : 1;
	28562 : 1;
	28563 : 1;
	28564 : 1;
	28565 : 1;
	28566 : 1;
	28567 : 1;
	28568 : 1;
	28569 : 1;
	28570 : 1;
	28571 : 1;
	28572 : 1;
	28573 : 1;
	28574 : 1;
	28575 : 1;
	28576 : 1;
	28577 : 1;
	28578 : 1;
	28579 : 1;
	28580 : 1;
	28581 : 1;
	28582 : 1;
	28583 : 1;
	28584 : 1;
	28585 : 1;
	28586 : 1;
	28587 : 1;
	28588 : 1;
	28589 : 1;
	28590 : 1;
	28591 : 1;
	28592 : 1;
	28593 : 1;
	28594 : 1;
	28595 : 1;
	28596 : 1;
	28597 : 1;
	28598 : 0;
	28599 : 0;
	28600 : 0;
	28601 : 1;
	28602 : 1;
	28603 : 1;
	28604 : 1;
	28605 : 1;
	28606 : 1;
	28607 : 1;
	28608 : 1;
	28609 : 1;
	28610 : 1;
	28611 : 1;
	28612 : 1;
	28613 : 1;
	28614 : 1;
	28615 : 1;
	28616 : 1;
	28617 : 1;
	28618 : 1;
	28619 : 1;
	28620 : 1;
	28621 : 1;
	28622 : 1;
	28623 : 1;
	28624 : 1;
	28625 : 1;
	28626 : 1;
	28627 : 1;
	28628 : 1;
	28629 : 1;
	28630 : 1;
	28631 : 1;
	28632 : 1;
	28633 : 1;
	28634 : 1;
	28635 : 1;
	28636 : 0;
	28637 : 0;
	28638 : 0;
	28639 : 0;
	28640 : 0;
	28641 : 1;
	28642 : 1;
	28643 : 1;
	28644 : 1;
	28645 : 1;
	28646 : 1;
	28647 : 1;
	28648 : 1;
	28649 : 1;
	28650 : 1;
	28651 : 1;
	28652 : 1;
	28653 : 1;
	28654 : 1;
	28655 : 1;
	28656 : 1;
	28657 : 1;
	28658 : 1;
	28659 : 1;
	28660 : 1;
	28661 : 1;
	28662 : 1;
	28663 : 1;
	28664 : 1;
	28665 : 1;
	28666 : 1;
	28667 : 1;
	28668 : 1;
	28669 : 1;
	28670 : 1;
	28671 : 1;
	28672 : 1;
	28673 : 0;
	28674 : 0;
	28675 : 0;
	28676 : 1;
	28677 : 1;
	28678 : 1;
	28679 : 1;
	28680 : 1;
	28681 : 1;
	28682 : 1;
	28683 : 1;
	28684 : 1;
	28685 : 1;
	28686 : 1;
	28687 : 1;
	28688 : 1;
	28689 : 1;
	28690 : 1;
	28691 : 1;
	28692 : 1;
	28693 : 1;
	28694 : 1;
	28695 : 1;
	28696 : 1;
	28697 : 1;
	28698 : 1;
	28699 : 1;
	28700 : 1;
	28701 : 1;
	28702 : 1;
	28703 : 1;
	28704 : 1;
	28705 : 1;
	28706 : 1;
	28707 : 1;
	28708 : 1;
	28709 : 1;
	28710 : 1;
	28711 : 1;
	28712 : 1;
	28713 : 1;
	28714 : 1;
	28715 : 1;
	28716 : 1;
	28717 : 1;
	28718 : 1;
	28719 : 1;
	28720 : 1;
	28721 : 1;
	28722 : 0;
	28723 : 0;
	28724 : 0;
	28725 : 1;
	28726 : 1;
	28727 : 0;
	28728 : 1;
	28729 : 1;
	28730 : 1;
	28731 : 1;
	28732 : 1;
	28733 : 1;
	28734 : 1;
	28735 : 1;
	28736 : 1;
	28737 : 1;
	28738 : 1;
	28739 : 1;
	28740 : 1;
	28741 : 1;
	28742 : 1;
	28743 : 1;
	28744 : 1;
	28745 : 1;
	28746 : 1;
	28747 : 1;
	28748 : 1;
	28749 : 1;
	28750 : 1;
	28751 : 1;
	28752 : 1;
	28753 : 1;
	28754 : 1;
	28755 : 1;
	28756 : 1;
	28757 : 1;
	28758 : 1;
	28759 : 1;
	28760 : 1;
	28761 : 1;
	28762 : 1;
	28763 : 1;
	28764 : 1;
	28765 : 1;
	28766 : 1;
	28767 : 1;
	28768 : 1;
	28769 : 1;
	28770 : 1;
	28771 : 1;
	28772 : 1;
	28773 : 1;
	28774 : 1;
	28775 : 1;
	28776 : 1;
	28777 : 1;
	28778 : 1;
	28779 : 1;
	28780 : 1;
	28781 : 1;
	28782 : 1;
	28783 : 1;
	28784 : 1;
	28785 : 1;
	28786 : 1;
	28787 : 1;
	28788 : 1;
	28789 : 1;
	28790 : 1;
	28791 : 1;
	28792 : 1;
	28793 : 1;
	28794 : 1;
	28795 : 1;
	28796 : 1;
	28797 : 1;
	28798 : 1;
	28799 : 1;
	28800 : 1;
	28801 : 1;
	28802 : 1;
	28803 : 1;
	28804 : 1;
	28805 : 1;
	28806 : 1;
	28807 : 1;
	28808 : 1;
	28809 : 1;
	28810 : 1;
	28811 : 1;
	28812 : 1;
	28813 : 1;
	28814 : 1;
	28815 : 1;
	28816 : 1;
	28817 : 1;
	28818 : 1;
	28819 : 1;
	28820 : 1;
	28821 : 1;
	28822 : 1;
	28823 : 1;
	28824 : 1;
	28825 : 1;
	28826 : 1;
	28827 : 1;
	28828 : 1;
	28829 : 1;
	28830 : 1;
	28831 : 1;
	28832 : 1;
	28833 : 1;
	28834 : 1;
	28835 : 1;
	28836 : 1;
	28837 : 1;
	28838 : 1;
	28839 : 1;
	28840 : 1;
	28841 : 1;
	28842 : 1;
	28843 : 1;
	28844 : 1;
	28845 : 1;
	28846 : 1;
	28847 : 1;
	28848 : 1;
	28849 : 1;
	28850 : 1;
	28851 : 1;
	28852 : 1;
	28853 : 1;
	28854 : 1;
	28855 : 1;
	28856 : 1;
	28857 : 1;
	28858 : 1;
	28859 : 1;
	28860 : 1;
	28861 : 1;
	28862 : 1;
	28863 : 1;
	28864 : 1;
	28865 : 1;
	28866 : 1;
	28867 : 1;
	28868 : 1;
	28869 : 1;
	28870 : 1;
	28871 : 1;
	28872 : 1;
	28873 : 1;
	28874 : 1;
	28875 : 1;
	28876 : 1;
	28877 : 1;
	28878 : 1;
	28879 : 1;
	28880 : 1;
	28881 : 1;
	28882 : 1;
	28883 : 1;
	28884 : 1;
	28885 : 1;
	28886 : 1;
	28887 : 1;
	28888 : 1;
	28889 : 1;
	28890 : 1;
	28891 : 1;
	28892 : 1;
	28893 : 1;
	28894 : 1;
	28895 : 1;
	28896 : 1;
	28897 : 1;
	28898 : 1;
	28899 : 1;
	28900 : 1;
	28901 : 1;
	28902 : 1;
	28903 : 1;
	28904 : 1;
	28905 : 1;
	28906 : 1;
	28907 : 1;
	28908 : 1;
	28909 : 1;
	28910 : 1;
	28911 : 1;
	28912 : 1;
	28913 : 1;
	28914 : 1;
	28915 : 1;
	28916 : 1;
	28917 : 1;
	28918 : 1;
	28919 : 1;
	28920 : 1;
	28921 : 1;
	28922 : 1;
	28923 : 1;
	28924 : 1;
	28925 : 1;
	28926 : 1;
	28927 : 1;
	28928 : 1;
	28929 : 1;
	28930 : 1;
	28931 : 1;
	28932 : 1;
	28933 : 1;
	28934 : 1;
	28935 : 1;
	28936 : 1;
	28937 : 1;
	28938 : 1;
	28939 : 1;
	28940 : 1;
	28941 : 1;
	28942 : 1;
	28943 : 1;
	28944 : 1;
	28945 : 1;
	28946 : 1;
	28947 : 1;
	28948 : 1;
	28949 : 1;
	28950 : 1;
	28951 : 1;
	28952 : 1;
	28953 : 1;
	28954 : 1;
	28955 : 1;
	28956 : 1;
	28957 : 1;
	28958 : 1;
	28959 : 1;
	28960 : 1;
	28961 : 1;
	28962 : 1;
	28963 : 1;
	28964 : 1;
	28965 : 1;
	28966 : 1;
	28967 : 1;
	28968 : 1;
	28969 : 1;
	28970 : 1;
	28971 : 1;
	28972 : 1;
	28973 : 1;
	28974 : 1;
	28975 : 1;
	28976 : 1;
	28977 : 1;
	28978 : 1;
	28979 : 1;
	28980 : 1;
	28981 : 1;
	28982 : 1;
	28983 : 1;
	28984 : 1;
	28985 : 1;
	28986 : 1;
	28987 : 1;
	28988 : 1;
	28989 : 1;
	28990 : 1;
	28991 : 1;
	28992 : 1;
	28993 : 1;
	28994 : 1;
	28995 : 1;
	28996 : 1;
	28997 : 1;
	28998 : 1;
	28999 : 1;
	29000 : 1;
	29001 : 1;
	29002 : 1;
	29003 : 1;
	29004 : 1;
	29005 : 1;
	29006 : 1;
	29007 : 1;
	29008 : 1;
	29009 : 1;
	29010 : 1;
	29011 : 1;
	29012 : 1;
	29013 : 1;
	29014 : 1;
	29015 : 1;
	29016 : 1;
	29017 : 1;
	29018 : 1;
	29019 : 1;
	29020 : 1;
	29021 : 1;
	29022 : 1;
	29023 : 1;
	29024 : 1;
	29025 : 1;
	29026 : 1;
	29027 : 1;
	29028 : 1;
	29029 : 1;
	29030 : 1;
	29031 : 1;
	29032 : 1;
	29033 : 1;
	29034 : 1;
	29035 : 1;
	29036 : 1;
	29037 : 1;
	29038 : 1;
	29039 : 1;
	29040 : 1;
	29041 : 1;
	29042 : 1;
	29043 : 1;
	29044 : 1;
	29045 : 1;
	29046 : 1;
	29047 : 1;
	29048 : 1;
	29049 : 1;
	29050 : 1;
	29051 : 1;
	29052 : 1;
	29053 : 1;
	29054 : 1;
	29055 : 1;
	29056 : 1;
	29057 : 1;
	29058 : 1;
	29059 : 1;
	29060 : 1;
	29061 : 1;
	29062 : 1;
	29063 : 1;
	29064 : 1;
	29065 : 1;
	29066 : 1;
	29067 : 1;
	29068 : 1;
	29069 : 1;
	29070 : 1;
	29071 : 1;
	29072 : 1;
	29073 : 1;
	29074 : 1;
	29075 : 1;
	29076 : 1;
	29077 : 1;
	29078 : 1;
	29079 : 1;
	29080 : 1;
	29081 : 1;
	29082 : 1;
	29083 : 1;
	29084 : 1;
	29085 : 1;
	29086 : 1;
	29087 : 1;
	29088 : 1;
	29089 : 1;
	29090 : 1;
	29091 : 1;
	29092 : 1;
	29093 : 1;
	29094 : 1;
	29095 : 1;
	29096 : 1;
	29097 : 1;
	29098 : 1;
	29099 : 1;
	29100 : 1;
	29101 : 1;
	29102 : 1;
	29103 : 1;
	29104 : 1;
	29105 : 1;
	29106 : 1;
	29107 : 1;
	29108 : 1;
	29109 : 1;
	29110 : 1;
	29111 : 1;
	29112 : 1;
	29113 : 1;
	29114 : 1;
	29115 : 1;
	29116 : 1;
	29117 : 1;
	29118 : 1;
	29119 : 1;
	29120 : 1;
	29121 : 1;
	29122 : 1;
	29123 : 1;
	29124 : 1;
	29125 : 1;
	29126 : 1;
	29127 : 1;
	29128 : 1;
	29129 : 1;
	29130 : 1;
	29131 : 1;
	29132 : 1;
	29133 : 1;
	29134 : 1;
	29135 : 1;
	29136 : 1;
	29137 : 1;
	29138 : 1;
	29139 : 1;
	29140 : 1;
	29141 : 1;
	29142 : 1;
	29143 : 1;
	29144 : 1;
	29145 : 1;
	29146 : 1;
	29147 : 1;
	29148 : 1;
	29149 : 1;
	29150 : 1;
	29151 : 1;
	29152 : 1;
	29153 : 1;
	29154 : 1;
	29155 : 1;
	29156 : 1;
	29157 : 1;
	29158 : 1;
	29159 : 1;
	29160 : 1;
	29161 : 1;
	29162 : 1;
	29163 : 1;
	29164 : 1;
	29165 : 1;
	29166 : 1;
	29167 : 1;
	29168 : 1;
	29169 : 1;
	29170 : 1;
	29171 : 1;
	29172 : 1;
	29173 : 1;
	29174 : 1;
	29175 : 1;
	29176 : 1;
	29177 : 1;
	29178 : 1;
	29179 : 1;
	29180 : 1;
	29181 : 1;
	29182 : 1;
	29183 : 1;
	29184 : 1;
	29185 : 1;
	29186 : 1;
	29187 : 1;
	29188 : 1;
	29189 : 1;
	29190 : 1;
	29191 : 1;
	29192 : 1;
	29193 : 1;
	29194 : 1;
	29195 : 1;
	29196 : 1;
	29197 : 1;
	29198 : 1;
	29199 : 1;
	29200 : 1;
	29201 : 1;
	29202 : 1;
	29203 : 1;
	29204 : 1;
	29205 : 1;
	29206 : 1;
	29207 : 1;
	29208 : 1;
	29209 : 1;
	29210 : 1;
	29211 : 1;
	29212 : 1;
	29213 : 1;
	29214 : 1;
	29215 : 1;
	29216 : 1;
	29217 : 1;
	29218 : 1;
	29219 : 1;
	29220 : 1;
	29221 : 1;
	29222 : 1;
	29223 : 1;
	29224 : 1;
	29225 : 1;
	29226 : 1;
	29227 : 1;
	29228 : 1;
	29229 : 1;
	29230 : 1;
	29231 : 1;
	29232 : 1;
	29233 : 1;
	29234 : 1;
	29235 : 1;
	29236 : 1;
	29237 : 1;
	29238 : 1;
	29239 : 1;
	29240 : 1;
	29241 : 1;
	29242 : 1;
	29243 : 1;
	29244 : 1;
	29245 : 1;
	29246 : 1;
	29247 : 1;
	29248 : 1;
	29249 : 1;
	29250 : 1;
	29251 : 1;
	29252 : 1;
	29253 : 1;
	29254 : 1;
	29255 : 1;
	29256 : 1;
	29257 : 1;
	29258 : 1;
	29259 : 1;
	29260 : 1;
	29261 : 1;
	29262 : 1;
	29263 : 1;
	29264 : 1;
	29265 : 1;
	29266 : 1;
	29267 : 1;
	29268 : 1;
	29269 : 1;
	29270 : 1;
	29271 : 1;
	29272 : 1;
	29273 : 1;
	29274 : 1;
	29275 : 1;
	29276 : 1;
	29277 : 1;
	29278 : 1;
	29279 : 1;
	29280 : 1;
	29281 : 1;
	29282 : 1;
	29283 : 1;
	29284 : 1;
	29285 : 1;
	29286 : 1;
	29287 : 1;
	29288 : 1;
	29289 : 1;
	29290 : 1;
	29291 : 1;
	29292 : 1;
	29293 : 1;
	29294 : 1;
	29295 : 1;
	29296 : 1;
	29297 : 1;
	29298 : 1;
	29299 : 1;
	29300 : 1;
	29301 : 1;
	29302 : 1;
	29303 : 1;
	29304 : 1;
	29305 : 1;
	29306 : 1;
	29307 : 1;
	29308 : 1;
	29309 : 1;
	29310 : 1;
	29311 : 1;
	29312 : 1;
	29313 : 1;
	29314 : 1;
	29315 : 1;
	29316 : 1;
	29317 : 1;
	29318 : 1;
	29319 : 1;
	29320 : 1;
	29321 : 1;
	29322 : 1;
	29323 : 1;
	29324 : 1;
	29325 : 1;
	29326 : 1;
	29327 : 1;
	29328 : 1;
	29329 : 1;
	29330 : 1;
	29331 : 1;
	29332 : 1;
	29333 : 1;
	29334 : 1;
	29335 : 1;
	29336 : 1;
	29337 : 1;
	29338 : 1;
	29339 : 1;
	29340 : 1;
	29341 : 1;
	29342 : 1;
	29343 : 1;
	29344 : 1;
	29345 : 1;
	29346 : 1;
	29347 : 1;
	29348 : 1;
	29349 : 1;
	29350 : 1;
	29351 : 1;
	29352 : 1;
	29353 : 1;
	29354 : 1;
	29355 : 1;
	29356 : 1;
	29357 : 1;
	29358 : 1;
	29359 : 1;
	29360 : 1;
	29361 : 1;
	29362 : 1;
	29363 : 1;
	29364 : 1;
	29365 : 1;
	29366 : 1;
	29367 : 1;
	29368 : 1;
	29369 : 1;
	29370 : 1;
	29371 : 1;
	29372 : 1;
	29373 : 1;
	29374 : 1;
	29375 : 1;
	29376 : 1;
	29377 : 1;
	29378 : 1;
	29379 : 1;
	29380 : 1;
	29381 : 1;
	29382 : 1;
	29383 : 1;
	29384 : 1;
	29385 : 1;
	29386 : 1;
	29387 : 1;
	29388 : 1;
	29389 : 1;
	29390 : 1;
	29391 : 1;
	29392 : 1;
	29393 : 1;
	29394 : 1;
	29395 : 1;
	29396 : 1;
	29397 : 1;
	29398 : 1;
	29399 : 1;
	29400 : 1;
	29401 : 1;
	29402 : 1;
	29403 : 1;
	29404 : 1;
	29405 : 1;
	29406 : 1;
	29407 : 1;
	29408 : 1;
	29409 : 1;
	29410 : 1;
	29411 : 1;
	29412 : 1;
	29413 : 1;
	29414 : 1;
	29415 : 1;
	29416 : 1;
	29417 : 1;
	29418 : 1;
	29419 : 1;
	29420 : 1;
	29421 : 1;
	29422 : 1;
	29423 : 1;
	29424 : 1;
	29425 : 1;
	29426 : 1;
	29427 : 1;
	29428 : 1;
	29429 : 1;
	29430 : 1;
	29431 : 1;
	29432 : 1;
	29433 : 1;
	29434 : 1;
	29435 : 1;
	29436 : 1;
	29437 : 1;
	29438 : 1;
	29439 : 1;
	29440 : 1;
	29441 : 1;
	29442 : 1;
	29443 : 1;
	29444 : 1;
	29445 : 1;
	29446 : 1;
	29447 : 1;
	29448 : 1;
	29449 : 1;
	29450 : 1;
	29451 : 1;
	29452 : 1;
	29453 : 1;
	29454 : 1;
	29455 : 1;
	29456 : 1;
	29457 : 1;
	29458 : 1;
	29459 : 1;
	29460 : 1;
	29461 : 1;
	29462 : 1;
	29463 : 1;
	29464 : 1;
	29465 : 1;
	29466 : 1;
	29467 : 1;
	29468 : 1;
	29469 : 1;
	29470 : 1;
	29471 : 1;
	29472 : 1;
	29473 : 1;
	29474 : 1;
	29475 : 1;
	29476 : 1;
	29477 : 1;
	29478 : 1;
	29479 : 1;
	29480 : 1;
	29481 : 1;
	29482 : 1;
	29483 : 1;
	29484 : 1;
	29485 : 1;
	29486 : 1;
	29487 : 1;
	29488 : 1;
	29489 : 1;
	29490 : 1;
	29491 : 1;
	29492 : 1;
	29493 : 1;
	29494 : 1;
	29495 : 1;
	29496 : 1;
	29497 : 1;
	29498 : 1;
	29499 : 1;
	29500 : 1;
	29501 : 1;
	29502 : 1;
	29503 : 1;
	29504 : 1;
	29505 : 1;
	29506 : 1;
	29507 : 1;
	29508 : 1;
	29509 : 1;
	29510 : 1;
	29511 : 1;
	29512 : 1;
	29513 : 1;
	29514 : 1;
	29515 : 1;
	29516 : 1;
	29517 : 1;
	29518 : 1;
	29519 : 1;
	29520 : 1;
	29521 : 1;
	29522 : 1;
	29523 : 1;
	29524 : 1;
	29525 : 1;
	29526 : 1;
	29527 : 1;
	29528 : 1;
	29529 : 1;
	29530 : 1;
	29531 : 1;
	29532 : 1;
	29533 : 1;
	29534 : 1;
	29535 : 1;
	29536 : 1;
	29537 : 1;
	29538 : 1;
	29539 : 1;
	29540 : 1;
	29541 : 1;
	29542 : 1;
	29543 : 1;
	29544 : 1;
	29545 : 1;
	29546 : 1;
	29547 : 1;
	29548 : 1;
	29549 : 1;
	29550 : 1;
	29551 : 1;
	29552 : 1;
	29553 : 1;
	29554 : 1;
	29555 : 1;
	29556 : 1;
	29557 : 1;
	29558 : 1;
	29559 : 1;
	29560 : 1;
	29561 : 1;
	29562 : 1;
	29563 : 1;
	29564 : 1;
	29565 : 1;
	29566 : 1;
	29567 : 1;
	29568 : 1;
	29569 : 1;
	29570 : 1;
	29571 : 1;
	29572 : 1;
	29573 : 1;
	29574 : 1;
	29575 : 1;
	29576 : 1;
	29577 : 1;
	29578 : 1;
	29579 : 1;
	29580 : 1;
	29581 : 1;
	29582 : 1;
	29583 : 1;
	29584 : 1;
	29585 : 1;
	29586 : 1;
	29587 : 1;
	29588 : 1;
	29589 : 1;
	29590 : 1;
	29591 : 1;
	29592 : 1;
	29593 : 1;
	29594 : 1;
	29595 : 1;
	29596 : 1;
	29597 : 1;
	29598 : 1;
	29599 : 1;
	29600 : 1;
	29601 : 1;
	29602 : 1;
	29603 : 1;
	29604 : 1;
	29605 : 1;
	29606 : 1;
	29607 : 1;
	29608 : 1;
	29609 : 1;
	29610 : 1;
	29611 : 1;
	29612 : 1;
	29613 : 1;
	29614 : 1;
	29615 : 1;
	29616 : 1;
	29617 : 1;
	29618 : 1;
	29619 : 1;
	29620 : 1;
	29621 : 1;
	29622 : 1;
	29623 : 1;
	29624 : 1;
	29625 : 1;
	29626 : 1;
	29627 : 1;
	29628 : 1;
	29629 : 1;
	29630 : 1;
	29631 : 1;
	29632 : 1;
	29633 : 1;
	29634 : 1;
	29635 : 1;
	29636 : 1;
	29637 : 1;
	29638 : 1;
	29639 : 1;
	29640 : 1;
	29641 : 1;
	29642 : 1;
	29643 : 1;
	29644 : 1;
	29645 : 1;
	29646 : 1;
	29647 : 1;
	29648 : 1;
	29649 : 1;
	29650 : 1;
	29651 : 1;
	29652 : 1;
	29653 : 1;
	29654 : 1;
	29655 : 1;
	29656 : 1;
	29657 : 1;
	29658 : 1;
	29659 : 1;
	29660 : 1;
	29661 : 1;
	29662 : 1;
	29663 : 1;
	29664 : 1;
	29665 : 1;
	29666 : 1;
	29667 : 1;
	29668 : 1;
	29669 : 1;
	29670 : 1;
	29671 : 1;
	29672 : 1;
	29673 : 1;
	29674 : 1;
	29675 : 1;
	29676 : 1;
	29677 : 1;
	29678 : 1;
	29679 : 1;
	29680 : 1;
	29681 : 1;
	29682 : 1;
	29683 : 1;
	29684 : 1;
	29685 : 1;
	29686 : 1;
	29687 : 1;
	29688 : 1;
	29689 : 1;
	29690 : 1;
	29691 : 1;
	29692 : 1;
	29693 : 1;
	29694 : 1;
	29695 : 1;
	29696 : 1;
	29697 : 1;
	29698 : 1;
	29699 : 1;
	29700 : 1;
	29701 : 1;
	29702 : 1;
	29703 : 1;
	29704 : 1;
	29705 : 1;
	29706 : 1;
	29707 : 1;
	29708 : 1;
	29709 : 1;
	29710 : 1;
	29711 : 1;
	29712 : 1;
	29713 : 1;
	29714 : 1;
	29715 : 1;
	29716 : 1;
	29717 : 1;
	29718 : 1;
	29719 : 1;
	29720 : 1;
	29721 : 1;
	29722 : 1;
	29723 : 1;
	29724 : 1;
	29725 : 1;
	29726 : 1;
	29727 : 1;
	29728 : 1;
	29729 : 1;
	29730 : 1;
	29731 : 1;
	29732 : 1;
	29733 : 1;
	29734 : 1;
	29735 : 1;
	29736 : 1;
	29737 : 1;
	29738 : 1;
	29739 : 1;
	29740 : 1;
	29741 : 1;
	29742 : 1;
	29743 : 1;
	29744 : 1;
	29745 : 1;
	29746 : 1;
	29747 : 1;
	29748 : 1;
	29749 : 1;
	29750 : 1;
	29751 : 1;
	29752 : 1;
	29753 : 1;
	29754 : 1;
	29755 : 1;
	29756 : 1;
	29757 : 1;
	29758 : 1;
	29759 : 1;
	29760 : 1;
	29761 : 1;
	29762 : 1;
	29763 : 1;
	29764 : 1;
	29765 : 1;
	29766 : 1;
	29767 : 1;
	29768 : 1;
	29769 : 1;
	29770 : 1;
	29771 : 1;
	29772 : 1;
	29773 : 1;
	29774 : 1;
	29775 : 1;
	29776 : 1;
	29777 : 1;
	29778 : 1;
	29779 : 1;
	29780 : 1;
	29781 : 1;
	29782 : 1;
	29783 : 1;
	29784 : 1;
	29785 : 1;
	29786 : 1;
	29787 : 1;
	29788 : 1;
	29789 : 1;
	29790 : 1;
	29791 : 1;
	29792 : 1;
	29793 : 1;
	29794 : 1;
	29795 : 1;
	29796 : 1;
	29797 : 1;
	29798 : 1;
	29799 : 1;
	29800 : 1;
	29801 : 1;
	29802 : 1;
	29803 : 1;
	29804 : 1;
	29805 : 1;
	29806 : 1;
	29807 : 1;
	29808 : 1;
	29809 : 1;
	29810 : 1;
	29811 : 1;
	29812 : 1;
	29813 : 1;
	29814 : 1;
	29815 : 1;
	29816 : 1;
	29817 : 1;
	29818 : 1;
	29819 : 1;
	29820 : 1;
	29821 : 1;
	29822 : 1;
	29823 : 1;
	29824 : 1;
	29825 : 1;
	29826 : 1;
	29827 : 1;
	29828 : 1;
	29829 : 1;
	29830 : 1;
	29831 : 1;
	29832 : 1;
	29833 : 1;
	29834 : 1;
	29835 : 1;
	29836 : 1;
	29837 : 1;
	29838 : 1;
	29839 : 1;
	29840 : 1;
	29841 : 1;
	29842 : 1;
	29843 : 1;
	29844 : 1;
	29845 : 1;
	29846 : 1;
	29847 : 1;
	29848 : 1;
	29849 : 1;
	29850 : 1;
	29851 : 1;
	29852 : 1;
	29853 : 1;
	29854 : 1;
	29855 : 1;
	29856 : 1;
	29857 : 1;
	29858 : 1;
	29859 : 1;
	29860 : 1;
	29861 : 1;
	29862 : 1;
	29863 : 1;
	29864 : 1;
	29865 : 1;
	29866 : 1;
	29867 : 1;
	29868 : 1;
	29869 : 1;
	29870 : 1;
	29871 : 1;
	29872 : 1;
	29873 : 1;
	29874 : 1;
	29875 : 1;
	29876 : 1;
	29877 : 1;
	29878 : 1;
	29879 : 1;
	29880 : 1;
	29881 : 1;
	29882 : 1;
	29883 : 1;
	29884 : 1;
	29885 : 1;
	29886 : 1;
	29887 : 1;
	29888 : 1;
	29889 : 1;
	29890 : 1;
	29891 : 1;
	29892 : 1;
	29893 : 1;
	29894 : 1;
	29895 : 1;
	29896 : 1;
	29897 : 1;
	29898 : 1;
	29899 : 1;
	29900 : 1;
	29901 : 1;
	29902 : 1;
	29903 : 1;
	29904 : 1;
	29905 : 1;
	29906 : 1;
	29907 : 1;
	29908 : 1;
	29909 : 1;
	29910 : 1;
	29911 : 1;
	29912 : 1;
	29913 : 1;
	29914 : 1;
	29915 : 1;
	29916 : 1;
	29917 : 1;
	29918 : 1;
	29919 : 1;
	29920 : 1;
	29921 : 1;
	29922 : 1;
	29923 : 1;
	29924 : 1;
	29925 : 1;
	29926 : 1;
	29927 : 1;
	29928 : 1;
	29929 : 1;
	29930 : 1;
	29931 : 1;
	29932 : 1;
	29933 : 1;
	29934 : 1;
	29935 : 1;
	29936 : 1;
	29937 : 1;
	29938 : 1;
	29939 : 1;
	29940 : 1;
	29941 : 1;
	29942 : 1;
	29943 : 1;
	29944 : 1;
	29945 : 1;
	29946 : 1;
	29947 : 1;
	29948 : 1;
	29949 : 1;
	29950 : 1;
	29951 : 1;
	29952 : 1;
	29953 : 1;
	29954 : 1;
	29955 : 1;
	29956 : 1;
	29957 : 1;
	29958 : 1;
	29959 : 1;
	29960 : 1;
	29961 : 1;
	29962 : 1;
	29963 : 1;
	29964 : 1;
	29965 : 1;
	29966 : 1;
	29967 : 1;
	29968 : 1;
	29969 : 1;
	29970 : 1;
	29971 : 1;
	29972 : 1;
	29973 : 1;
	29974 : 1;
	29975 : 1;
	29976 : 1;
	29977 : 1;
	29978 : 1;
	29979 : 1;
	29980 : 1;
	29981 : 1;
	29982 : 1;
	29983 : 1;
	29984 : 1;
	29985 : 1;
	29986 : 1;
	29987 : 1;
	29988 : 1;
	29989 : 1;
	29990 : 1;
	29991 : 1;
	29992 : 1;
	29993 : 1;
	29994 : 1;
	29995 : 1;
	29996 : 1;
	29997 : 1;
	29998 : 1;
	29999 : 1;
	30000 : 1;
	30001 : 1;
	30002 : 1;
	30003 : 1;
	30004 : 1;
	30005 : 1;
	30006 : 1;
	30007 : 1;
	30008 : 1;
	30009 : 1;
	30010 : 1;
	30011 : 1;
	30012 : 1;
	30013 : 1;
	30014 : 1;
	30015 : 1;
	30016 : 1;
	30017 : 1;
	30018 : 1;
	30019 : 1;
	30020 : 1;
	30021 : 1;
	30022 : 1;
	30023 : 1;
	30024 : 1;
	30025 : 1;
	30026 : 1;
	30027 : 1;
	30028 : 1;
	30029 : 1;
	30030 : 1;
	30031 : 1;
	30032 : 1;
	30033 : 1;
	30034 : 1;
	30035 : 1;
	30036 : 1;
	30037 : 1;
	30038 : 1;
	30039 : 1;
	30040 : 1;
	30041 : 1;
	30042 : 1;
	30043 : 1;
	30044 : 1;
	30045 : 1;
	30046 : 1;
	30047 : 1;
	30048 : 1;
	30049 : 1;
	30050 : 1;
	30051 : 1;
	30052 : 1;
	30053 : 1;
	30054 : 1;
	30055 : 1;
	30056 : 1;
	30057 : 1;
	30058 : 1;
	30059 : 1;
	30060 : 1;
	30061 : 1;
	30062 : 1;
	30063 : 1;
	30064 : 1;
	30065 : 1;
	30066 : 1;
	30067 : 1;
	30068 : 1;
	30069 : 1;
	30070 : 1;
	30071 : 1;
	30072 : 1;
	30073 : 1;
	30074 : 1;
	30075 : 1;
	30076 : 1;
	30077 : 1;
	30078 : 1;
	30079 : 1;
	30080 : 1;
	30081 : 1;
	30082 : 1;
	30083 : 1;
	30084 : 1;
	30085 : 1;
	30086 : 1;
	30087 : 1;
	30088 : 1;
	30089 : 1;
	30090 : 1;
	30091 : 1;
	30092 : 1;
	30093 : 1;
	30094 : 1;
	30095 : 1;
	30096 : 1;
	30097 : 1;
	30098 : 1;
	30099 : 1;
	30100 : 1;
	30101 : 1;
	30102 : 1;
	30103 : 1;
	30104 : 1;
	30105 : 1;
	30106 : 1;
	30107 : 1;
	30108 : 1;
	30109 : 1;
	30110 : 1;
	30111 : 1;
	30112 : 1;
	30113 : 1;
	30114 : 1;
	30115 : 1;
	30116 : 1;
	30117 : 1;
	30118 : 1;
	30119 : 1;
	30120 : 1;
	30121 : 1;
	30122 : 1;
	30123 : 1;
	30124 : 1;
	30125 : 1;
	30126 : 1;
	30127 : 1;
	30128 : 1;
	30129 : 1;
	30130 : 1;
	30131 : 1;
	30132 : 1;
	30133 : 1;
	30134 : 1;
	30135 : 1;
	30136 : 1;
	30137 : 1;
	30138 : 1;
	30139 : 1;
	30140 : 1;
	30141 : 1;
	30142 : 1;
	30143 : 1;
	30144 : 1;
	30145 : 1;
	30146 : 1;
	30147 : 1;
	30148 : 1;
	30149 : 1;
	30150 : 1;
	30151 : 1;
	30152 : 1;
	30153 : 1;
	30154 : 1;
	30155 : 1;
	30156 : 1;
	30157 : 1;
	30158 : 1;
	30159 : 1;
	30160 : 1;
	30161 : 1;
	30162 : 1;
	30163 : 1;
	30164 : 1;
	30165 : 1;
	30166 : 1;
	30167 : 1;
	30168 : 1;
	30169 : 1;
	30170 : 1;
	30171 : 1;
	30172 : 1;
	30173 : 1;
	30174 : 1;
	30175 : 1;
	30176 : 1;
	30177 : 1;
	30178 : 1;
	30179 : 1;
	30180 : 1;
	30181 : 1;
	30182 : 1;
	30183 : 1;
	30184 : 1;
	30185 : 1;
	30186 : 1;
	30187 : 1;
	30188 : 1;
	30189 : 1;
	30190 : 1;
	30191 : 1;
	30192 : 1;
	30193 : 1;
	30194 : 1;
	30195 : 1;
	30196 : 1;
	30197 : 1;
	30198 : 1;
	30199 : 1;
	30200 : 1;
	30201 : 1;
	30202 : 1;
	30203 : 1;
	30204 : 1;
	30205 : 1;
	30206 : 1;
	30207 : 1;
	30208 : 1;
	30209 : 1;
	30210 : 1;
	30211 : 1;
	30212 : 1;
	30213 : 1;
	30214 : 1;
	30215 : 1;
	30216 : 1;
	30217 : 1;
	30218 : 1;
	30219 : 1;
	30220 : 1;
	30221 : 1;
	30222 : 1;
	30223 : 1;
	30224 : 1;
	30225 : 1;
	30226 : 1;
	30227 : 1;
	30228 : 1;
	30229 : 1;
	30230 : 1;
	30231 : 1;
	30232 : 1;
	30233 : 1;
	30234 : 1;
	30235 : 1;
	30236 : 1;
	30237 : 1;
	30238 : 1;
	30239 : 1;
	30240 : 1;
	30241 : 1;
	30242 : 1;
	30243 : 1;
	30244 : 1;
	30245 : 1;
	30246 : 1;
	30247 : 1;
	30248 : 1;
	30249 : 1;
	30250 : 1;
	30251 : 1;
	30252 : 1;
	30253 : 1;
	30254 : 1;
	30255 : 1;
	30256 : 1;
	30257 : 1;
	30258 : 1;
	30259 : 1;
	30260 : 1;
	30261 : 1;
	30262 : 1;
	30263 : 1;
	30264 : 1;
	30265 : 1;
	30266 : 1;
	30267 : 1;
	30268 : 1;
	30269 : 1;
	30270 : 1;
	30271 : 1;
	30272 : 1;
	30273 : 1;
	30274 : 1;
	30275 : 1;
	30276 : 1;
	30277 : 1;
	30278 : 1;
	30279 : 1;
	30280 : 1;
	30281 : 1;
	30282 : 1;
	30283 : 1;
	30284 : 1;
	30285 : 1;
	30286 : 1;
	30287 : 1;
	30288 : 1;
	30289 : 1;
	30290 : 1;
	30291 : 1;
	30292 : 1;
	30293 : 1;
	30294 : 1;
	30295 : 1;
	30296 : 1;
	30297 : 1;
	30298 : 1;
	30299 : 1;
	30300 : 1;
	30301 : 1;
	30302 : 1;
	30303 : 1;
	30304 : 1;
	30305 : 1;
	30306 : 1;
	30307 : 1;
	30308 : 1;
	30309 : 1;
	30310 : 1;
	30311 : 1;
	30312 : 1;
	30313 : 1;
	30314 : 1;
	30315 : 1;
	30316 : 1;
	30317 : 1;
	30318 : 1;
	30319 : 1;
	30320 : 1;
	30321 : 1;
	30322 : 1;
	30323 : 1;
	30324 : 1;
	30325 : 1;
	30326 : 1;
	30327 : 1;
	30328 : 1;
	30329 : 1;
	30330 : 1;
	30331 : 1;
	30332 : 1;
	30333 : 1;
	30334 : 1;
	30335 : 1;
	30336 : 1;
	30337 : 1;
	30338 : 1;
	30339 : 1;
	30340 : 1;
	30341 : 1;
	30342 : 1;
	30343 : 1;
	30344 : 1;
	30345 : 1;
	30346 : 1;
	30347 : 1;
	30348 : 1;
	30349 : 1;
	30350 : 1;
	30351 : 1;
	30352 : 1;
	30353 : 1;
	30354 : 1;
	30355 : 1;
	30356 : 1;
	30357 : 1;
	30358 : 1;
	30359 : 1;
	30360 : 1;
	30361 : 1;
	30362 : 1;
	30363 : 1;
	30364 : 1;
	30365 : 1;
	30366 : 1;
	30367 : 1;
	30368 : 1;
	30369 : 1;
	30370 : 1;
	30371 : 1;
	30372 : 1;
	30373 : 1;
	30374 : 1;
	30375 : 1;
	30376 : 1;
	30377 : 1;
	30378 : 1;
	30379 : 1;
	30380 : 1;
	30381 : 1;
	30382 : 1;
	30383 : 1;
	30384 : 1;
	30385 : 1;
	30386 : 1;
	30387 : 1;
	30388 : 1;
	30389 : 1;
	30390 : 1;
	30391 : 1;
	30392 : 1;
	30393 : 1;
	30394 : 1;
	30395 : 1;
	30396 : 1;
	30397 : 1;
	30398 : 1;
	30399 : 1;
	30400 : 1;
	30401 : 1;
	30402 : 1;
	30403 : 1;
	30404 : 1;
	30405 : 1;
	30406 : 1;
	30407 : 1;
	30408 : 1;
	30409 : 1;
	30410 : 1;
	30411 : 1;
	30412 : 1;
	30413 : 1;
	30414 : 1;
	30415 : 1;
	30416 : 1;
	30417 : 1;
	30418 : 1;
	30419 : 1;
	30420 : 1;
	30421 : 1;
	30422 : 1;
	30423 : 1;
	30424 : 1;
	30425 : 1;
	30426 : 1;
	30427 : 1;
	30428 : 1;
	30429 : 1;
	30430 : 1;
	30431 : 1;
	30432 : 1;
	30433 : 1;
	30434 : 1;
	30435 : 1;
	30436 : 1;
	30437 : 1;
	30438 : 1;
	30439 : 1;
	30440 : 1;
	30441 : 1;
	30442 : 1;
	30443 : 1;
	30444 : 1;
	30445 : 1;
	30446 : 1;
	30447 : 1;
	30448 : 1;
	30449 : 1;
	30450 : 1;
	30451 : 1;
	30452 : 1;
	30453 : 1;
	30454 : 1;
	30455 : 1;
	30456 : 1;
	30457 : 1;
	30458 : 1;
	30459 : 1;
	30460 : 1;
	30461 : 1;
	30462 : 1;
	30463 : 1;
	30464 : 1;
	30465 : 1;
	30466 : 1;
	30467 : 1;
	30468 : 1;
	30469 : 1;
	30470 : 1;
	30471 : 1;
	30472 : 1;
	30473 : 1;
	30474 : 1;
	30475 : 1;
	30476 : 1;
	30477 : 1;
	30478 : 1;
	30479 : 1;
	30480 : 1;
	30481 : 1;
	30482 : 1;
	30483 : 1;
	30484 : 1;
	30485 : 1;
	30486 : 1;
	30487 : 1;
	30488 : 1;
	30489 : 1;
	30490 : 1;
	30491 : 1;
	30492 : 1;
	30493 : 1;
	30494 : 1;
	30495 : 1;
	30496 : 1;
	30497 : 1;
	30498 : 1;
	30499 : 1;
	30500 : 1;
	30501 : 1;
	30502 : 1;
	30503 : 1;
	30504 : 1;
	30505 : 1;
	30506 : 1;
	30507 : 1;
	30508 : 1;
	30509 : 1;
	30510 : 1;
	30511 : 1;
	30512 : 1;
	30513 : 1;
	30514 : 1;
	30515 : 1;
	30516 : 1;
	30517 : 1;
	30518 : 1;
	30519 : 1;
	30520 : 1;
	30521 : 1;
	30522 : 1;
	30523 : 1;
	30524 : 1;
	30525 : 1;
	30526 : 1;
	30527 : 1;
	30528 : 1;
	30529 : 1;
	30530 : 1;
	30531 : 1;
	30532 : 1;
	30533 : 1;
	30534 : 1;
	30535 : 1;
	30536 : 1;
	30537 : 1;
	30538 : 1;
	30539 : 1;
	30540 : 1;
	30541 : 1;
	30542 : 1;
	30543 : 1;
	30544 : 1;
	30545 : 1;
	30546 : 1;
	30547 : 1;
	30548 : 1;
	30549 : 1;
	30550 : 1;
	30551 : 1;
	30552 : 1;
	30553 : 1;
	30554 : 1;
	30555 : 1;
	30556 : 1;
	30557 : 1;
	30558 : 1;
	30559 : 1;
	30560 : 1;
	30561 : 1;
	30562 : 1;
	30563 : 1;
	30564 : 1;
	30565 : 1;
	30566 : 1;
	30567 : 1;
	30568 : 1;
	30569 : 1;
	30570 : 1;
	30571 : 1;
	30572 : 1;
	30573 : 1;
	30574 : 1;
	30575 : 1;
	30576 : 1;
	30577 : 1;
	30578 : 1;
	30579 : 1;
	30580 : 1;
	30581 : 1;
	30582 : 1;
	30583 : 1;
	30584 : 1;
	30585 : 1;
	30586 : 1;
	30587 : 1;
	30588 : 1;
	30589 : 1;
	30590 : 1;
	30591 : 1;
	30592 : 1;
	30593 : 1;
	30594 : 1;
	30595 : 1;
	30596 : 1;
	30597 : 1;
	30598 : 1;
	30599 : 1;
	30600 : 1;
	30601 : 1;
	30602 : 1;
	30603 : 1;
	30604 : 1;
	30605 : 1;
	30606 : 1;
	30607 : 1;
	30608 : 1;
	30609 : 1;
	30610 : 1;
	30611 : 1;
	30612 : 1;
	30613 : 1;
	30614 : 1;
	30615 : 1;
	30616 : 1;
	30617 : 1;
	30618 : 1;
	30619 : 1;
	30620 : 1;
	30621 : 1;
	30622 : 1;
	30623 : 1;
	30624 : 1;
	30625 : 1;
	30626 : 1;
	30627 : 1;
	30628 : 1;
	30629 : 1;
	30630 : 1;
	30631 : 1;
	30632 : 1;
	30633 : 1;
	30634 : 1;
	30635 : 1;
	30636 : 1;
	30637 : 1;
	30638 : 1;
	30639 : 1;
	30640 : 1;
	30641 : 1;
	30642 : 1;
	30643 : 1;
	30644 : 1;
	30645 : 1;
	30646 : 1;
	30647 : 1;
	30648 : 1;
	30649 : 1;
	30650 : 1;
	30651 : 1;
	30652 : 1;
	30653 : 1;
	30654 : 1;
	30655 : 1;
	30656 : 1;
	30657 : 1;
	30658 : 1;
	30659 : 1;
	30660 : 1;
	30661 : 1;
	30662 : 1;
	30663 : 1;
	30664 : 1;
	30665 : 1;
	30666 : 1;
	30667 : 1;
	30668 : 1;
	30669 : 1;
	30670 : 1;
	30671 : 1;
	30672 : 1;
	30673 : 1;
	30674 : 1;
	30675 : 1;
	30676 : 1;
	30677 : 1;
	30678 : 1;
	30679 : 1;
	30680 : 1;
	30681 : 1;
	30682 : 1;
	30683 : 1;
	30684 : 1;
	30685 : 1;
	30686 : 1;
	30687 : 1;
	30688 : 1;
	30689 : 1;
	30690 : 1;
	30691 : 1;
	30692 : 1;
	30693 : 1;
	30694 : 1;
	30695 : 1;
	30696 : 1;
	30697 : 1;
	30698 : 1;
	30699 : 1;
	30700 : 1;
	30701 : 1;
	30702 : 1;
	30703 : 1;
	30704 : 1;
	30705 : 1;
	30706 : 1;
	30707 : 1;
	30708 : 1;
	30709 : 1;
	30710 : 1;
	30711 : 1;
	30712 : 1;
	30713 : 1;
	30714 : 1;
	30715 : 1;
	30716 : 1;
	30717 : 1;
	30718 : 1;
	30719 : 1;
	30720 : 1;
	30721 : 1;
	30722 : 1;
	30723 : 1;
	30724 : 1;
	30725 : 1;
	30726 : 1;
	30727 : 1;
	30728 : 1;
	30729 : 1;
	30730 : 1;
	30731 : 1;
	30732 : 1;
	30733 : 1;
	30734 : 1;
	30735 : 1;
	30736 : 1;
	30737 : 1;
	30738 : 1;
	30739 : 1;
	30740 : 1;
	30741 : 1;
	30742 : 1;
	30743 : 1;
	30744 : 1;
	30745 : 1;
	30746 : 1;
	30747 : 1;
	30748 : 1;
	30749 : 1;
	30750 : 1;
	30751 : 1;
	30752 : 1;
	30753 : 1;
	30754 : 1;
	30755 : 1;
	30756 : 1;
	30757 : 1;
	30758 : 1;
	30759 : 1;
	30760 : 1;
	30761 : 1;
	30762 : 1;
	30763 : 1;
	30764 : 1;
	30765 : 1;
	30766 : 1;
	30767 : 1;
	30768 : 1;
	30769 : 1;
	30770 : 1;
	30771 : 1;
	30772 : 1;
	30773 : 1;
	30774 : 1;
	30775 : 1;
	30776 : 1;
	30777 : 1;
	30778 : 1;
	30779 : 1;
	30780 : 1;
	30781 : 1;
	30782 : 1;
	30783 : 1;
	30784 : 1;
	30785 : 1;
	30786 : 1;
	30787 : 1;
	30788 : 1;
	30789 : 1;
	30790 : 1;
	30791 : 1;
	30792 : 1;
	30793 : 1;
	30794 : 1;
	30795 : 1;
	30796 : 1;
	30797 : 1;
	30798 : 1;
	30799 : 1;
	30800 : 1;
	30801 : 1;
	30802 : 1;
	30803 : 1;
	30804 : 1;
	30805 : 1;
	30806 : 1;
	30807 : 1;
	30808 : 1;
	30809 : 1;
	30810 : 1;
	30811 : 1;
	30812 : 1;
	30813 : 1;
	30814 : 1;
	30815 : 1;
	30816 : 1;
	30817 : 1;
	30818 : 1;
	30819 : 1;
	30820 : 1;
	30821 : 1;
	30822 : 1;
	30823 : 1;
	30824 : 1;
	30825 : 1;
	30826 : 1;
	30827 : 1;
	30828 : 1;
	30829 : 1;
	30830 : 1;
	30831 : 1;
	30832 : 1;
	30833 : 1;
	30834 : 1;
	30835 : 1;
	30836 : 0;
	30837 : 0;
	30838 : 1;
	30839 : 1;
	30840 : 1;
	30841 : 1;
	30842 : 1;
	30843 : 1;
	30844 : 1;
	30845 : 1;
	30846 : 1;
	30847 : 1;
	30848 : 1;
	30849 : 1;
	30850 : 1;
	30851 : 1;
	30852 : 1;
	30853 : 1;
	30854 : 1;
	30855 : 1;
	30856 : 1;
	30857 : 1;
	30858 : 1;
	30859 : 1;
	30860 : 1;
	30861 : 1;
	30862 : 1;
	30863 : 1;
	30864 : 1;
	30865 : 1;
	30866 : 1;
	30867 : 1;
	30868 : 1;
	30869 : 1;
	30870 : 1;
	30871 : 1;
	30872 : 1;
	30873 : 1;
	30874 : 1;
	30875 : 1;
	30876 : 1;
	30877 : 1;
	30878 : 1;
	30879 : 1;
	30880 : 1;
	30881 : 1;
	30882 : 1;
	30883 : 1;
	30884 : 1;
	30885 : 1;
	30886 : 1;
	30887 : 1;
	30888 : 1;
	30889 : 1;
	30890 : 1;
	30891 : 1;
	30892 : 1;
	30893 : 1;
	30894 : 1;
	30895 : 1;
	30896 : 1;
	30897 : 1;
	30898 : 1;
	30899 : 1;
	30900 : 1;
	30901 : 1;
	30902 : 1;
	30903 : 1;
	30904 : 1;
	30905 : 1;
	30906 : 1;
	30907 : 1;
	30908 : 1;
	30909 : 1;
	30910 : 1;
	30911 : 1;
	30912 : 1;
	30913 : 1;
	30914 : 1;
	30915 : 1;
	30916 : 1;
	30917 : 1;
	30918 : 1;
	30919 : 1;
	30920 : 1;
	30921 : 1;
	30922 : 1;
	30923 : 1;
	30924 : 1;
	30925 : 1;
	30926 : 1;
	30927 : 1;
	30928 : 1;
	30929 : 1;
	30930 : 1;
	30931 : 1;
	30932 : 1;
	30933 : 1;
	30934 : 1;
	30935 : 1;
	30936 : 1;
	30937 : 1;
	30938 : 1;
	30939 : 1;
	30940 : 1;
	30941 : 1;
	30942 : 1;
	30943 : 1;
	30944 : 1;
	30945 : 1;
	30946 : 1;
	30947 : 1;
	30948 : 1;
	30949 : 1;
	30950 : 1;
	30951 : 1;
	30952 : 1;
	30953 : 1;
	30954 : 1;
	30955 : 1;
	30956 : 1;
	30957 : 1;
	30958 : 1;
	30959 : 1;
	30960 : 1;
	30961 : 1;
	30962 : 1;
	30963 : 1;
	30964 : 1;
	30965 : 1;
	30966 : 1;
	30967 : 1;
	30968 : 1;
	30969 : 1;
	30970 : 1;
	30971 : 1;
	30972 : 1;
	30973 : 1;
	30974 : 1;
	30975 : 1;
	30976 : 1;
	30977 : 1;
	30978 : 1;
	30979 : 1;
	30980 : 1;
	30981 : 1;
	30982 : 1;
	30983 : 1;
	30984 : 1;
	30985 : 1;
	30986 : 1;
	30987 : 1;
	30988 : 1;
	30989 : 1;
	30990 : 1;
	30991 : 1;
	30992 : 1;
	30993 : 1;
	30994 : 1;
	30995 : 1;
	30996 : 1;
	30997 : 1;
	30998 : 1;
	30999 : 1;
	31000 : 1;
	31001 : 1;
	31002 : 1;
	31003 : 1;
	31004 : 1;
	31005 : 1;
	31006 : 1;
	31007 : 1;
	31008 : 1;
	31009 : 1;
	31010 : 1;
	31011 : 1;
	31012 : 1;
	31013 : 1;
	31014 : 1;
	31015 : 1;
	31016 : 1;
	31017 : 1;
	31018 : 1;
	31019 : 1;
	31020 : 1;
	31021 : 1;
	31022 : 1;
	31023 : 1;
	31024 : 1;
	31025 : 1;
	31026 : 1;
	31027 : 1;
	31028 : 1;
	31029 : 1;
	31030 : 1;
	31031 : 1;
	31032 : 1;
	31033 : 1;
	31034 : 1;
	31035 : 1;
	31036 : 1;
	31037 : 1;
	31038 : 1;
	31039 : 1;
	31040 : 1;
	31041 : 1;
	31042 : 1;
	31043 : 1;
	31044 : 1;
	31045 : 1;
	31046 : 1;
	31047 : 1;
	31048 : 1;
	31049 : 1;
	31050 : 1;
	31051 : 1;
	31052 : 1;
	31053 : 1;
	31054 : 1;
	31055 : 1;
	31056 : 1;
	31057 : 1;
	31058 : 1;
	31059 : 1;
	31060 : 1;
	31061 : 1;
	31062 : 1;
	31063 : 1;
	31064 : 1;
	31065 : 1;
	31066 : 1;
	31067 : 1;
	31068 : 1;
	31069 : 1;
	31070 : 1;
	31071 : 1;
	31072 : 1;
	31073 : 1;
	31074 : 1;
	31075 : 1;
	31076 : 0;
	31077 : 0;
	31078 : 1;
	31079 : 1;
	31080 : 1;
	31081 : 1;
	31082 : 1;
	31083 : 1;
	31084 : 1;
	31085 : 1;
	31086 : 1;
	31087 : 1;
	31088 : 1;
	31089 : 1;
	31090 : 1;
	31091 : 1;
	31092 : 1;
	31093 : 1;
	31094 : 1;
	31095 : 1;
	31096 : 1;
	31097 : 1;
	31098 : 1;
	31099 : 1;
	31100 : 1;
	31101 : 1;
	31102 : 1;
	31103 : 1;
	31104 : 1;
	31105 : 1;
	31106 : 1;
	31107 : 1;
	31108 : 1;
	31109 : 1;
	31110 : 1;
	31111 : 1;
	31112 : 1;
	31113 : 1;
	31114 : 1;
	31115 : 1;
	31116 : 1;
	31117 : 1;
	31118 : 1;
	31119 : 1;
	31120 : 1;
	31121 : 1;
	31122 : 1;
	31123 : 1;
	31124 : 1;
	31125 : 1;
	31126 : 1;
	31127 : 1;
	31128 : 1;
	31129 : 1;
	31130 : 1;
	31131 : 1;
	31132 : 1;
	31133 : 1;
	31134 : 1;
	31135 : 1;
	31136 : 1;
	31137 : 1;
	31138 : 1;
	31139 : 1;
	31140 : 1;
	31141 : 1;
	31142 : 1;
	31143 : 1;
	31144 : 1;
	31145 : 1;
	31146 : 1;
	31147 : 1;
	31148 : 1;
	31149 : 1;
	31150 : 1;
	31151 : 1;
	31152 : 1;
	31153 : 1;
	31154 : 1;
	31155 : 1;
	31156 : 1;
	31157 : 1;
	31158 : 1;
	31159 : 1;
	31160 : 1;
	31161 : 1;
	31162 : 1;
	31163 : 1;
	31164 : 1;
	31165 : 1;
	31166 : 1;
	31167 : 1;
	31168 : 1;
	31169 : 1;
	31170 : 1;
	31171 : 1;
	31172 : 1;
	31173 : 1;
	31174 : 1;
	31175 : 1;
	31176 : 1;
	31177 : 1;
	31178 : 1;
	31179 : 1;
	31180 : 1;
	31181 : 1;
	31182 : 1;
	31183 : 1;
	31184 : 1;
	31185 : 1;
	31186 : 1;
	31187 : 1;
	31188 : 1;
	31189 : 1;
	31190 : 1;
	31191 : 1;
	31192 : 1;
	31193 : 1;
	31194 : 1;
	31195 : 1;
	31196 : 1;
	31197 : 1;
	31198 : 1;
	31199 : 1;
	31200 : 1;
	31201 : 1;
	31202 : 1;
	31203 : 1;
	31204 : 1;
	31205 : 1;
	31206 : 1;
	31207 : 1;
	31208 : 1;
	31209 : 1;
	31210 : 1;
	31211 : 1;
	31212 : 1;
	31213 : 1;
	31214 : 1;
	31215 : 1;
	31216 : 1;
	31217 : 1;
	31218 : 1;
	31219 : 1;
	31220 : 1;
	31221 : 1;
	31222 : 1;
	31223 : 1;
	31224 : 1;
	31225 : 1;
	31226 : 1;
	31227 : 1;
	31228 : 1;
	31229 : 1;
	31230 : 1;
	31231 : 1;
	31232 : 1;
	31233 : 1;
	31234 : 1;
	31235 : 1;
	31236 : 1;
	31237 : 1;
	31238 : 1;
	31239 : 1;
	31240 : 1;
	31241 : 1;
	31242 : 1;
	31243 : 1;
	31244 : 1;
	31245 : 1;
	31246 : 1;
	31247 : 1;
	31248 : 1;
	31249 : 1;
	31250 : 1;
	31251 : 1;
	31252 : 1;
	31253 : 1;
	31254 : 1;
	31255 : 1;
	31256 : 1;
	31257 : 1;
	31258 : 1;
	31259 : 1;
	31260 : 1;
	31261 : 1;
	31262 : 1;
	31263 : 1;
	31264 : 1;
	31265 : 1;
	31266 : 1;
	31267 : 1;
	31268 : 1;
	31269 : 1;
	31270 : 1;
	31271 : 1;
	31272 : 1;
	31273 : 1;
	31274 : 1;
	31275 : 1;
	31276 : 1;
	31277 : 1;
	31278 : 1;
	31279 : 1;
	31280 : 1;
	31281 : 1;
	31282 : 1;
	31283 : 1;
	31284 : 1;
	31285 : 1;
	31286 : 1;
	31287 : 1;
	31288 : 1;
	31289 : 1;
	31290 : 1;
	31291 : 1;
	31292 : 1;
	31293 : 1;
	31294 : 1;
	31295 : 1;
	31296 : 1;
	31297 : 1;
	31298 : 1;
	31299 : 1;
	31300 : 1;
	31301 : 1;
	31302 : 1;
	31303 : 1;
	31304 : 1;
	31305 : 1;
	31306 : 1;
	31307 : 1;
	31308 : 1;
	31309 : 1;
	31310 : 1;
	31311 : 1;
	31312 : 1;
	31313 : 1;
	31314 : 1;
	31315 : 1;
	31316 : 0;
	31317 : 0;
	31318 : 1;
	31319 : 1;
	31320 : 1;
	31321 : 1;
	31322 : 1;
	31323 : 1;
	31324 : 1;
	31325 : 1;
	31326 : 1;
	31327 : 1;
	31328 : 1;
	31329 : 1;
	31330 : 0;
	31331 : 0;
	31332 : 0;
	31333 : 0;
	31334 : 1;
	31335 : 1;
	31336 : 1;
	31337 : 1;
	31338 : 1;
	31339 : 1;
	31340 : 1;
	31341 : 1;
	31342 : 1;
	31343 : 1;
	31344 : 1;
	31345 : 1;
	31346 : 1;
	31347 : 1;
	31348 : 1;
	31349 : 1;
	31350 : 1;
	31351 : 1;
	31352 : 1;
	31353 : 1;
	31354 : 1;
	31355 : 1;
	31356 : 1;
	31357 : 1;
	31358 : 1;
	31359 : 1;
	31360 : 1;
	31361 : 1;
	31362 : 1;
	31363 : 1;
	31364 : 1;
	31365 : 1;
	31366 : 1;
	31367 : 1;
	31368 : 1;
	31369 : 1;
	31370 : 1;
	31371 : 0;
	31372 : 1;
	31373 : 1;
	31374 : 1;
	31375 : 0;
	31376 : 0;
	31377 : 0;
	31378 : 0;
	31379 : 0;
	31380 : 1;
	31381 : 1;
	31382 : 1;
	31383 : 1;
	31384 : 1;
	31385 : 1;
	31386 : 1;
	31387 : 0;
	31388 : 1;
	31389 : 0;
	31390 : 0;
	31391 : 1;
	31392 : 1;
	31393 : 1;
	31394 : 1;
	31395 : 1;
	31396 : 1;
	31397 : 1;
	31398 : 1;
	31399 : 1;
	31400 : 1;
	31401 : 1;
	31402 : 1;
	31403 : 1;
	31404 : 1;
	31405 : 1;
	31406 : 1;
	31407 : 1;
	31408 : 1;
	31409 : 1;
	31410 : 1;
	31411 : 1;
	31412 : 1;
	31413 : 1;
	31414 : 1;
	31415 : 1;
	31416 : 1;
	31417 : 1;
	31418 : 1;
	31419 : 1;
	31420 : 1;
	31421 : 1;
	31422 : 1;
	31423 : 1;
	31424 : 1;
	31425 : 1;
	31426 : 1;
	31427 : 1;
	31428 : 1;
	31429 : 1;
	31430 : 1;
	31431 : 1;
	31432 : 1;
	31433 : 1;
	31434 : 1;
	31435 : 1;
	31436 : 1;
	31437 : 1;
	31438 : 1;
	31439 : 1;
	31440 : 1;
	31441 : 1;
	31442 : 1;
	31443 : 1;
	31444 : 1;
	31445 : 1;
	31446 : 1;
	31447 : 1;
	31448 : 1;
	31449 : 1;
	31450 : 1;
	31451 : 1;
	31452 : 1;
	31453 : 1;
	31454 : 1;
	31455 : 1;
	31456 : 1;
	31457 : 1;
	31458 : 1;
	31459 : 1;
	31460 : 1;
	31461 : 1;
	31462 : 1;
	31463 : 1;
	31464 : 1;
	31465 : 1;
	31466 : 1;
	31467 : 1;
	31468 : 1;
	31469 : 1;
	31470 : 1;
	31471 : 1;
	31472 : 1;
	31473 : 1;
	31474 : 1;
	31475 : 1;
	31476 : 1;
	31477 : 1;
	31478 : 1;
	31479 : 1;
	31480 : 1;
	31481 : 1;
	31482 : 1;
	31483 : 1;
	31484 : 1;
	31485 : 1;
	31486 : 1;
	31487 : 1;
	31488 : 1;
	31489 : 1;
	31490 : 1;
	31491 : 1;
	31492 : 1;
	31493 : 1;
	31494 : 1;
	31495 : 1;
	31496 : 1;
	31497 : 1;
	31498 : 1;
	31499 : 1;
	31500 : 1;
	31501 : 1;
	31502 : 1;
	31503 : 1;
	31504 : 1;
	31505 : 1;
	31506 : 1;
	31507 : 1;
	31508 : 1;
	31509 : 1;
	31510 : 1;
	31511 : 1;
	31512 : 1;
	31513 : 1;
	31514 : 1;
	31515 : 0;
	31516 : 1;
	31517 : 1;
	31518 : 1;
	31519 : 1;
	31520 : 1;
	31521 : 1;
	31522 : 1;
	31523 : 1;
	31524 : 1;
	31525 : 1;
	31526 : 1;
	31527 : 1;
	31528 : 1;
	31529 : 1;
	31530 : 1;
	31531 : 1;
	31532 : 1;
	31533 : 1;
	31534 : 1;
	31535 : 1;
	31536 : 1;
	31537 : 1;
	31538 : 1;
	31539 : 1;
	31540 : 1;
	31541 : 1;
	31542 : 1;
	31543 : 1;
	31544 : 1;
	31545 : 1;
	31546 : 1;
	31547 : 1;
	31548 : 1;
	31549 : 1;
	31550 : 1;
	31551 : 1;
	31552 : 1;
	31553 : 1;
	31554 : 1;
	31555 : 1;
	31556 : 0;
	31557 : 0;
	31558 : 1;
	31559 : 1;
	31560 : 1;
	31561 : 1;
	31562 : 1;
	31563 : 1;
	31564 : 1;
	31565 : 1;
	31566 : 1;
	31567 : 1;
	31568 : 1;
	31569 : 0;
	31570 : 1;
	31571 : 1;
	31572 : 1;
	31573 : 0;
	31574 : 1;
	31575 : 1;
	31576 : 1;
	31577 : 1;
	31578 : 1;
	31579 : 1;
	31580 : 1;
	31581 : 1;
	31582 : 1;
	31583 : 1;
	31584 : 1;
	31585 : 1;
	31586 : 1;
	31587 : 1;
	31588 : 1;
	31589 : 1;
	31590 : 1;
	31591 : 1;
	31592 : 1;
	31593 : 1;
	31594 : 1;
	31595 : 1;
	31596 : 1;
	31597 : 1;
	31598 : 1;
	31599 : 1;
	31600 : 1;
	31601 : 1;
	31602 : 1;
	31603 : 1;
	31604 : 1;
	31605 : 1;
	31606 : 1;
	31607 : 1;
	31608 : 1;
	31609 : 1;
	31610 : 1;
	31611 : 0;
	31612 : 1;
	31613 : 1;
	31614 : 1;
	31615 : 0;
	31616 : 1;
	31617 : 1;
	31618 : 1;
	31619 : 1;
	31620 : 1;
	31621 : 1;
	31622 : 1;
	31623 : 1;
	31624 : 1;
	31625 : 1;
	31626 : 1;
	31627 : 1;
	31628 : 1;
	31629 : 1;
	31630 : 0;
	31631 : 1;
	31632 : 1;
	31633 : 1;
	31634 : 1;
	31635 : 1;
	31636 : 1;
	31637 : 1;
	31638 : 1;
	31639 : 1;
	31640 : 1;
	31641 : 1;
	31642 : 1;
	31643 : 1;
	31644 : 1;
	31645 : 1;
	31646 : 1;
	31647 : 1;
	31648 : 1;
	31649 : 1;
	31650 : 1;
	31651 : 1;
	31652 : 1;
	31653 : 1;
	31654 : 1;
	31655 : 1;
	31656 : 1;
	31657 : 1;
	31658 : 1;
	31659 : 1;
	31660 : 1;
	31661 : 1;
	31662 : 1;
	31663 : 1;
	31664 : 1;
	31665 : 1;
	31666 : 1;
	31667 : 1;
	31668 : 1;
	31669 : 1;
	31670 : 1;
	31671 : 1;
	31672 : 1;
	31673 : 1;
	31674 : 1;
	31675 : 1;
	31676 : 1;
	31677 : 1;
	31678 : 1;
	31679 : 1;
	31680 : 1;
	31681 : 1;
	31682 : 1;
	31683 : 1;
	31684 : 1;
	31685 : 1;
	31686 : 1;
	31687 : 1;
	31688 : 1;
	31689 : 1;
	31690 : 1;
	31691 : 1;
	31692 : 1;
	31693 : 1;
	31694 : 1;
	31695 : 1;
	31696 : 1;
	31697 : 1;
	31698 : 1;
	31699 : 1;
	31700 : 1;
	31701 : 1;
	31702 : 1;
	31703 : 1;
	31704 : 1;
	31705 : 1;
	31706 : 1;
	31707 : 1;
	31708 : 1;
	31709 : 1;
	31710 : 1;
	31711 : 1;
	31712 : 1;
	31713 : 1;
	31714 : 1;
	31715 : 1;
	31716 : 1;
	31717 : 1;
	31718 : 1;
	31719 : 1;
	31720 : 1;
	31721 : 1;
	31722 : 1;
	31723 : 1;
	31724 : 1;
	31725 : 1;
	31726 : 1;
	31727 : 1;
	31728 : 1;
	31729 : 1;
	31730 : 1;
	31731 : 1;
	31732 : 1;
	31733 : 1;
	31734 : 1;
	31735 : 1;
	31736 : 1;
	31737 : 1;
	31738 : 1;
	31739 : 1;
	31740 : 1;
	31741 : 1;
	31742 : 1;
	31743 : 1;
	31744 : 1;
	31745 : 1;
	31746 : 1;
	31747 : 1;
	31748 : 1;
	31749 : 1;
	31750 : 1;
	31751 : 1;
	31752 : 1;
	31753 : 1;
	31754 : 0;
	31755 : 0;
	31756 : 1;
	31757 : 1;
	31758 : 1;
	31759 : 1;
	31760 : 1;
	31761 : 1;
	31762 : 1;
	31763 : 1;
	31764 : 1;
	31765 : 1;
	31766 : 1;
	31767 : 1;
	31768 : 1;
	31769 : 1;
	31770 : 1;
	31771 : 1;
	31772 : 1;
	31773 : 1;
	31774 : 1;
	31775 : 1;
	31776 : 1;
	31777 : 1;
	31778 : 1;
	31779 : 1;
	31780 : 1;
	31781 : 1;
	31782 : 1;
	31783 : 1;
	31784 : 1;
	31785 : 1;
	31786 : 1;
	31787 : 1;
	31788 : 1;
	31789 : 1;
	31790 : 1;
	31791 : 1;
	31792 : 1;
	31793 : 1;
	31794 : 1;
	31795 : 1;
	31796 : 0;
	31797 : 0;
	31798 : 1;
	31799 : 1;
	31800 : 1;
	31801 : 1;
	31802 : 1;
	31803 : 1;
	31804 : 1;
	31805 : 1;
	31806 : 1;
	31807 : 1;
	31808 : 1;
	31809 : 0;
	31810 : 1;
	31811 : 1;
	31812 : 1;
	31813 : 0;
	31814 : 1;
	31815 : 1;
	31816 : 1;
	31817 : 1;
	31818 : 1;
	31819 : 1;
	31820 : 1;
	31821 : 1;
	31822 : 1;
	31823 : 1;
	31824 : 1;
	31825 : 1;
	31826 : 1;
	31827 : 1;
	31828 : 1;
	31829 : 1;
	31830 : 1;
	31831 : 1;
	31832 : 1;
	31833 : 1;
	31834 : 1;
	31835 : 1;
	31836 : 1;
	31837 : 1;
	31838 : 1;
	31839 : 1;
	31840 : 1;
	31841 : 1;
	31842 : 1;
	31843 : 1;
	31844 : 1;
	31845 : 1;
	31846 : 1;
	31847 : 1;
	31848 : 1;
	31849 : 1;
	31850 : 0;
	31851 : 0;
	31852 : 1;
	31853 : 1;
	31854 : 1;
	31855 : 0;
	31856 : 1;
	31857 : 1;
	31858 : 1;
	31859 : 1;
	31860 : 1;
	31861 : 1;
	31862 : 1;
	31863 : 1;
	31864 : 1;
	31865 : 1;
	31866 : 1;
	31867 : 1;
	31868 : 1;
	31869 : 1;
	31870 : 0;
	31871 : 1;
	31872 : 1;
	31873 : 1;
	31874 : 1;
	31875 : 1;
	31876 : 1;
	31877 : 1;
	31878 : 1;
	31879 : 1;
	31880 : 1;
	31881 : 1;
	31882 : 1;
	31883 : 1;
	31884 : 1;
	31885 : 1;
	31886 : 1;
	31887 : 1;
	31888 : 1;
	31889 : 1;
	31890 : 1;
	31891 : 1;
	31892 : 1;
	31893 : 1;
	31894 : 1;
	31895 : 1;
	31896 : 1;
	31897 : 1;
	31898 : 1;
	31899 : 1;
	31900 : 1;
	31901 : 1;
	31902 : 1;
	31903 : 1;
	31904 : 1;
	31905 : 1;
	31906 : 1;
	31907 : 1;
	31908 : 1;
	31909 : 1;
	31910 : 1;
	31911 : 1;
	31912 : 1;
	31913 : 1;
	31914 : 1;
	31915 : 1;
	31916 : 1;
	31917 : 1;
	31918 : 1;
	31919 : 1;
	31920 : 1;
	31921 : 1;
	31922 : 1;
	31923 : 1;
	31924 : 1;
	31925 : 1;
	31926 : 1;
	31927 : 1;
	31928 : 1;
	31929 : 1;
	31930 : 1;
	31931 : 1;
	31932 : 1;
	31933 : 1;
	31934 : 1;
	31935 : 1;
	31936 : 1;
	31937 : 1;
	31938 : 1;
	31939 : 1;
	31940 : 1;
	31941 : 1;
	31942 : 1;
	31943 : 1;
	31944 : 1;
	31945 : 1;
	31946 : 1;
	31947 : 1;
	31948 : 1;
	31949 : 1;
	31950 : 1;
	31951 : 1;
	31952 : 1;
	31953 : 1;
	31954 : 1;
	31955 : 1;
	31956 : 1;
	31957 : 1;
	31958 : 1;
	31959 : 1;
	31960 : 1;
	31961 : 1;
	31962 : 0;
	31963 : 0;
	31964 : 0;
	31965 : 0;
	31966 : 0;
	31967 : 1;
	31968 : 1;
	31969 : 1;
	31970 : 0;
	31971 : 0;
	31972 : 0;
	31973 : 0;
	31974 : 1;
	31975 : 1;
	31976 : 0;
	31977 : 1;
	31978 : 0;
	31979 : 0;
	31980 : 1;
	31981 : 1;
	31982 : 0;
	31983 : 0;
	31984 : 0;
	31985 : 0;
	31986 : 1;
	31987 : 1;
	31988 : 0;
	31989 : 0;
	31990 : 0;
	31991 : 0;
	31992 : 0;
	31993 : 1;
	31994 : 0;
	31995 : 0;
	31996 : 0;
	31997 : 0;
	31998 : 1;
	31999 : 1;
	32000 : 1;
	32001 : 0;
	32002 : 0;
	32003 : 0;
	32004 : 0;
	32005 : 1;
	32006 : 0;
	32007 : 1;
	32008 : 1;
	32009 : 0;
	32010 : 0;
	32011 : 1;
	32012 : 0;
	32013 : 0;
	32014 : 0;
	32015 : 0;
	32016 : 0;
	32017 : 1;
	32018 : 1;
	32019 : 0;
	32020 : 0;
	32021 : 0;
	32022 : 0;
	32023 : 1;
	32024 : 1;
	32025 : 1;
	32026 : 0;
	32027 : 0;
	32028 : 0;
	32029 : 0;
	32030 : 1;
	32031 : 0;
	32032 : 0;
	32033 : 0;
	32034 : 0;
	32035 : 1;
	32036 : 0;
	32037 : 0;
	32038 : 1;
	32039 : 1;
	32040 : 1;
	32041 : 1;
	32042 : 1;
	32043 : 0;
	32044 : 0;
	32045 : 0;
	32046 : 0;
	32047 : 0;
	32048 : 1;
	32049 : 0;
	32050 : 1;
	32051 : 1;
	32052 : 1;
	32053 : 0;
	32054 : 1;
	32055 : 0;
	32056 : 0;
	32057 : 0;
	32058 : 0;
	32059 : 1;
	32060 : 1;
	32061 : 0;
	32062 : 0;
	32063 : 0;
	32064 : 0;
	32065 : 1;
	32066 : 0;
	32067 : 0;
	32068 : 1;
	32069 : 1;
	32070 : 1;
	32071 : 0;
	32072 : 1;
	32073 : 1;
	32074 : 1;
	32075 : 1;
	32076 : 0;
	32077 : 0;
	32078 : 0;
	32079 : 0;
	32080 : 1;
	32081 : 0;
	32082 : 0;
	32083 : 0;
	32084 : 0;
	32085 : 1;
	32086 : 1;
	32087 : 0;
	32088 : 0;
	32089 : 0;
	32090 : 0;
	32091 : 0;
	32092 : 1;
	32093 : 1;
	32094 : 1;
	32095 : 0;
	32096 : 0;
	32097 : 0;
	32098 : 0;
	32099 : 1;
	32100 : 1;
	32101 : 0;
	32102 : 0;
	32103 : 0;
	32104 : 0;
	32105 : 0;
	32106 : 1;
	32107 : 0;
	32108 : 1;
	32109 : 1;
	32110 : 0;
	32111 : 1;
	32112 : 0;
	32113 : 0;
	32114 : 1;
	32115 : 1;
	32116 : 1;
	32117 : 0;
	32118 : 1;
	32119 : 1;
	32120 : 1;
	32121 : 1;
	32122 : 1;
	32123 : 1;
	32124 : 1;
	32125 : 1;
	32126 : 1;
	32127 : 1;
	32128 : 1;
	32129 : 1;
	32130 : 1;
	32131 : 1;
	32132 : 1;
	32133 : 1;
	32134 : 1;
	32135 : 1;
	32136 : 1;
	32137 : 1;
	32138 : 1;
	32139 : 1;
	32140 : 1;
	32141 : 1;
	32142 : 1;
	32143 : 1;
	32144 : 1;
	32145 : 1;
	32146 : 1;
	32147 : 1;
	32148 : 1;
	32149 : 1;
	32150 : 1;
	32151 : 1;
	32152 : 1;
	32153 : 1;
	32154 : 1;
	32155 : 1;
	32156 : 1;
	32157 : 1;
	32158 : 1;
	32159 : 1;
	32160 : 1;
	32161 : 1;
	32162 : 1;
	32163 : 1;
	32164 : 1;
	32165 : 1;
	32166 : 1;
	32167 : 1;
	32168 : 1;
	32169 : 1;
	32170 : 1;
	32171 : 1;
	32172 : 1;
	32173 : 1;
	32174 : 1;
	32175 : 1;
	32176 : 1;
	32177 : 1;
	32178 : 1;
	32179 : 1;
	32180 : 1;
	32181 : 1;
	32182 : 1;
	32183 : 1;
	32184 : 1;
	32185 : 1;
	32186 : 1;
	32187 : 1;
	32188 : 1;
	32189 : 1;
	32190 : 1;
	32191 : 1;
	32192 : 1;
	32193 : 1;
	32194 : 1;
	32195 : 1;
	32196 : 1;
	32197 : 1;
	32198 : 1;
	32199 : 1;
	32200 : 1;
	32201 : 0;
	32202 : 0;
	32203 : 1;
	32204 : 1;
	32205 : 1;
	32206 : 0;
	32207 : 1;
	32208 : 1;
	32209 : 1;
	32210 : 0;
	32211 : 1;
	32212 : 1;
	32213 : 1;
	32214 : 0;
	32215 : 1;
	32216 : 0;
	32217 : 0;
	32218 : 1;
	32219 : 1;
	32220 : 1;
	32221 : 0;
	32222 : 0;
	32223 : 1;
	32224 : 1;
	32225 : 0;
	32226 : 0;
	32227 : 0;
	32228 : 0;
	32229 : 1;
	32230 : 1;
	32231 : 1;
	32232 : 0;
	32233 : 1;
	32234 : 1;
	32235 : 0;
	32236 : 1;
	32237 : 1;
	32238 : 1;
	32239 : 1;
	32240 : 1;
	32241 : 0;
	32242 : 1;
	32243 : 1;
	32244 : 1;
	32245 : 1;
	32246 : 0;
	32247 : 1;
	32248 : 1;
	32249 : 0;
	32250 : 0;
	32251 : 1;
	32252 : 0;
	32253 : 0;
	32254 : 0;
	32255 : 0;
	32256 : 1;
	32257 : 0;
	32258 : 1;
	32259 : 0;
	32260 : 1;
	32261 : 0;
	32262 : 1;
	32263 : 0;
	32264 : 1;
	32265 : 0;
	32266 : 1;
	32267 : 1;
	32268 : 1;
	32269 : 0;
	32270 : 1;
	32271 : 0;
	32272 : 0;
	32273 : 1;
	32274 : 1;
	32275 : 1;
	32276 : 0;
	32277 : 0;
	32278 : 1;
	32279 : 1;
	32280 : 1;
	32281 : 1;
	32282 : 1;
	32283 : 1;
	32284 : 1;
	32285 : 1;
	32286 : 1;
	32287 : 1;
	32288 : 1;
	32289 : 0;
	32290 : 0;
	32291 : 0;
	32292 : 0;
	32293 : 0;
	32294 : 1;
	32295 : 0;
	32296 : 0;
	32297 : 1;
	32298 : 1;
	32299 : 1;
	32300 : 0;
	32301 : 1;
	32302 : 1;
	32303 : 1;
	32304 : 0;
	32305 : 0;
	32306 : 0;
	32307 : 0;
	32308 : 1;
	32309 : 1;
	32310 : 1;
	32311 : 0;
	32312 : 1;
	32313 : 1;
	32314 : 1;
	32315 : 0;
	32316 : 1;
	32317 : 1;
	32318 : 1;
	32319 : 0;
	32320 : 1;
	32321 : 0;
	32322 : 1;
	32323 : 1;
	32324 : 0;
	32325 : 0;
	32326 : 0;
	32327 : 0;
	32328 : 1;
	32329 : 1;
	32330 : 1;
	32331 : 0;
	32332 : 1;
	32333 : 1;
	32334 : 1;
	32335 : 0;
	32336 : 1;
	32337 : 1;
	32338 : 1;
	32339 : 1;
	32340 : 1;
	32341 : 0;
	32342 : 1;
	32343 : 0;
	32344 : 1;
	32345 : 0;
	32346 : 1;
	32347 : 0;
	32348 : 1;
	32349 : 1;
	32350 : 0;
	32351 : 1;
	32352 : 0;
	32353 : 0;
	32354 : 1;
	32355 : 1;
	32356 : 1;
	32357 : 0;
	32358 : 1;
	32359 : 1;
	32360 : 1;
	32361 : 1;
	32362 : 1;
	32363 : 1;
	32364 : 1;
	32365 : 1;
	32366 : 1;
	32367 : 1;
	32368 : 1;
	32369 : 1;
	32370 : 1;
	32371 : 1;
	32372 : 1;
	32373 : 1;
	32374 : 1;
	32375 : 1;
	32376 : 1;
	32377 : 1;
	32378 : 1;
	32379 : 1;
	32380 : 1;
	32381 : 1;
	32382 : 1;
	32383 : 1;
	32384 : 1;
	32385 : 1;
	32386 : 1;
	32387 : 1;
	32388 : 1;
	32389 : 1;
	32390 : 1;
	32391 : 1;
	32392 : 1;
	32393 : 1;
	32394 : 1;
	32395 : 1;
	32396 : 1;
	32397 : 1;
	32398 : 1;
	32399 : 1;
	32400 : 1;
	32401 : 1;
	32402 : 1;
	32403 : 1;
	32404 : 1;
	32405 : 1;
	32406 : 1;
	32407 : 1;
	32408 : 1;
	32409 : 1;
	32410 : 1;
	32411 : 1;
	32412 : 1;
	32413 : 1;
	32414 : 1;
	32415 : 1;
	32416 : 1;
	32417 : 1;
	32418 : 1;
	32419 : 1;
	32420 : 1;
	32421 : 1;
	32422 : 1;
	32423 : 1;
	32424 : 1;
	32425 : 1;
	32426 : 1;
	32427 : 1;
	32428 : 1;
	32429 : 1;
	32430 : 1;
	32431 : 1;
	32432 : 1;
	32433 : 1;
	32434 : 1;
	32435 : 1;
	32436 : 1;
	32437 : 1;
	32438 : 1;
	32439 : 1;
	32440 : 1;
	32441 : 0;
	32442 : 0;
	32443 : 1;
	32444 : 1;
	32445 : 1;
	32446 : 0;
	32447 : 1;
	32448 : 1;
	32449 : 1;
	32450 : 0;
	32451 : 1;
	32452 : 1;
	32453 : 1;
	32454 : 0;
	32455 : 1;
	32456 : 0;
	32457 : 1;
	32458 : 1;
	32459 : 1;
	32460 : 1;
	32461 : 0;
	32462 : 0;
	32463 : 0;
	32464 : 0;
	32465 : 0;
	32466 : 0;
	32467 : 0;
	32468 : 0;
	32469 : 1;
	32470 : 1;
	32471 : 1;
	32472 : 0;
	32473 : 1;
	32474 : 1;
	32475 : 0;
	32476 : 1;
	32477 : 1;
	32478 : 1;
	32479 : 1;
	32480 : 1;
	32481 : 1;
	32482 : 0;
	32483 : 0;
	32484 : 1;
	32485 : 1;
	32486 : 0;
	32487 : 1;
	32488 : 1;
	32489 : 0;
	32490 : 0;
	32491 : 1;
	32492 : 0;
	32493 : 0;
	32494 : 0;
	32495 : 0;
	32496 : 1;
	32497 : 0;
	32498 : 1;
	32499 : 0;
	32500 : 1;
	32501 : 0;
	32502 : 1;
	32503 : 0;
	32504 : 1;
	32505 : 0;
	32506 : 0;
	32507 : 0;
	32508 : 0;
	32509 : 0;
	32510 : 1;
	32511 : 0;
	32512 : 1;
	32513 : 1;
	32514 : 1;
	32515 : 1;
	32516 : 1;
	32517 : 1;
	32518 : 1;
	32519 : 1;
	32520 : 1;
	32521 : 1;
	32522 : 1;
	32523 : 1;
	32524 : 1;
	32525 : 1;
	32526 : 1;
	32527 : 1;
	32528 : 1;
	32529 : 0;
	32530 : 1;
	32531 : 1;
	32532 : 1;
	32533 : 0;
	32534 : 1;
	32535 : 0;
	32536 : 1;
	32537 : 1;
	32538 : 1;
	32539 : 1;
	32540 : 0;
	32541 : 1;
	32542 : 1;
	32543 : 1;
	32544 : 1;
	32545 : 1;
	32546 : 0;
	32547 : 0;
	32548 : 1;
	32549 : 1;
	32550 : 1;
	32551 : 0;
	32552 : 1;
	32553 : 1;
	32554 : 1;
	32555 : 0;
	32556 : 1;
	32557 : 1;
	32558 : 1;
	32559 : 0;
	32560 : 1;
	32561 : 0;
	32562 : 1;
	32563 : 1;
	32564 : 0;
	32565 : 0;
	32566 : 0;
	32567 : 0;
	32568 : 1;
	32569 : 1;
	32570 : 1;
	32571 : 0;
	32572 : 1;
	32573 : 1;
	32574 : 1;
	32575 : 0;
	32576 : 1;
	32577 : 1;
	32578 : 1;
	32579 : 1;
	32580 : 1;
	32581 : 0;
	32582 : 1;
	32583 : 0;
	32584 : 1;
	32585 : 0;
	32586 : 1;
	32587 : 0;
	32588 : 1;
	32589 : 1;
	32590 : 0;
	32591 : 1;
	32592 : 0;
	32593 : 0;
	32594 : 1;
	32595 : 1;
	32596 : 1;
	32597 : 0;
	32598 : 1;
	32599 : 1;
	32600 : 1;
	32601 : 1;
	32602 : 1;
	32603 : 1;
	32604 : 1;
	32605 : 1;
	32606 : 1;
	32607 : 1;
	32608 : 1;
	32609 : 1;
	32610 : 1;
	32611 : 1;
	32612 : 1;
	32613 : 1;
	32614 : 1;
	32615 : 1;
	32616 : 1;
	32617 : 1;
	32618 : 1;
	32619 : 1;
	32620 : 1;
	32621 : 1;
	32622 : 1;
	32623 : 1;
	32624 : 1;
	32625 : 1;
	32626 : 1;
	32627 : 1;
	32628 : 1;
	32629 : 1;
	32630 : 1;
	32631 : 1;
	32632 : 1;
	32633 : 1;
	32634 : 1;
	32635 : 1;
	32636 : 1;
	32637 : 1;
	32638 : 1;
	32639 : 1;
	32640 : 1;
	32641 : 1;
	32642 : 1;
	32643 : 1;
	32644 : 1;
	32645 : 1;
	32646 : 1;
	32647 : 1;
	32648 : 1;
	32649 : 1;
	32650 : 1;
	32651 : 1;
	32652 : 1;
	32653 : 1;
	32654 : 1;
	32655 : 1;
	32656 : 1;
	32657 : 1;
	32658 : 1;
	32659 : 1;
	32660 : 1;
	32661 : 1;
	32662 : 1;
	32663 : 1;
	32664 : 1;
	32665 : 1;
	32666 : 1;
	32667 : 1;
	32668 : 1;
	32669 : 1;
	32670 : 1;
	32671 : 1;
	32672 : 1;
	32673 : 1;
	32674 : 1;
	32675 : 1;
	32676 : 1;
	32677 : 1;
	32678 : 1;
	32679 : 1;
	32680 : 1;
	32681 : 0;
	32682 : 0;
	32683 : 1;
	32684 : 0;
	32685 : 0;
	32686 : 0;
	32687 : 1;
	32688 : 1;
	32689 : 1;
	32690 : 0;
	32691 : 1;
	32692 : 1;
	32693 : 1;
	32694 : 0;
	32695 : 1;
	32696 : 0;
	32697 : 1;
	32698 : 1;
	32699 : 1;
	32700 : 1;
	32701 : 0;
	32702 : 1;
	32703 : 1;
	32704 : 1;
	32705 : 1;
	32706 : 1;
	32707 : 0;
	32708 : 0;
	32709 : 1;
	32710 : 0;
	32711 : 0;
	32712 : 0;
	32713 : 1;
	32714 : 1;
	32715 : 0;
	32716 : 1;
	32717 : 1;
	32718 : 1;
	32719 : 1;
	32720 : 1;
	32721 : 1;
	32722 : 1;
	32723 : 1;
	32724 : 0;
	32725 : 1;
	32726 : 0;
	32727 : 1;
	32728 : 1;
	32729 : 0;
	32730 : 0;
	32731 : 1;
	32732 : 0;
	32733 : 0;
	32734 : 0;
	32735 : 0;
	32736 : 1;
	32737 : 0;
	32738 : 1;
	32739 : 0;
	32740 : 1;
	32741 : 0;
	32742 : 1;
	32743 : 0;
	32744 : 1;
	32745 : 0;
	32746 : 1;
	32747 : 1;
	32748 : 1;
	32749 : 1;
	32750 : 1;
	32751 : 0;
	32752 : 1;
	32753 : 1;
	32754 : 1;
	32755 : 1;
	32756 : 0;
	32757 : 0;
	32758 : 1;
	32759 : 1;
	32760 : 1;
	32761 : 1;
	32762 : 1;
	32763 : 1;
	32764 : 1;
	32765 : 1;
	32766 : 1;
	32767 : 1;
	32768 : 1;
	32769 : 0;
	32770 : 1;
	32771 : 1;
	32772 : 1;
	32773 : 0;
	32774 : 1;
	32775 : 0;
	32776 : 1;
	32777 : 1;
	32778 : 1;
	32779 : 1;
	32780 : 0;
	32781 : 1;
	32782 : 1;
	32783 : 1;
	32784 : 0;
	32785 : 0;
	32786 : 0;
	32787 : 0;
	32788 : 1;
	32789 : 1;
	32790 : 1;
	32791 : 0;
	32792 : 1;
	32793 : 1;
	32794 : 1;
	32795 : 0;
	32796 : 1;
	32797 : 1;
	32798 : 0;
	32799 : 0;
	32800 : 1;
	32801 : 0;
	32802 : 1;
	32803 : 1;
	32804 : 0;
	32805 : 0;
	32806 : 0;
	32807 : 0;
	32808 : 1;
	32809 : 1;
	32810 : 1;
	32811 : 0;
	32812 : 1;
	32813 : 1;
	32814 : 1;
	32815 : 0;
	32816 : 1;
	32817 : 1;
	32818 : 1;
	32819 : 1;
	32820 : 1;
	32821 : 0;
	32822 : 1;
	32823 : 0;
	32824 : 1;
	32825 : 0;
	32826 : 1;
	32827 : 0;
	32828 : 1;
	32829 : 1;
	32830 : 0;
	32831 : 1;
	32832 : 0;
	32833 : 0;
	32834 : 1;
	32835 : 1;
	32836 : 1;
	32837 : 0;
	32838 : 1;
	32839 : 1;
	32840 : 1;
	32841 : 1;
	32842 : 1;
	32843 : 1;
	32844 : 1;
	32845 : 1;
	32846 : 1;
	32847 : 1;
	32848 : 1;
	32849 : 1;
	32850 : 1;
	32851 : 1;
	32852 : 1;
	32853 : 1;
	32854 : 1;
	32855 : 1;
	32856 : 1;
	32857 : 1;
	32858 : 1;
	32859 : 1;
	32860 : 1;
	32861 : 1;
	32862 : 1;
	32863 : 1;
	32864 : 1;
	32865 : 1;
	32866 : 1;
	32867 : 1;
	32868 : 1;
	32869 : 1;
	32870 : 1;
	32871 : 1;
	32872 : 1;
	32873 : 1;
	32874 : 1;
	32875 : 1;
	32876 : 1;
	32877 : 1;
	32878 : 1;
	32879 : 1;
	32880 : 1;
	32881 : 1;
	32882 : 1;
	32883 : 1;
	32884 : 1;
	32885 : 1;
	32886 : 1;
	32887 : 1;
	32888 : 1;
	32889 : 1;
	32890 : 1;
	32891 : 1;
	32892 : 1;
	32893 : 1;
	32894 : 1;
	32895 : 1;
	32896 : 1;
	32897 : 1;
	32898 : 1;
	32899 : 1;
	32900 : 1;
	32901 : 1;
	32902 : 1;
	32903 : 1;
	32904 : 1;
	32905 : 1;
	32906 : 1;
	32907 : 1;
	32908 : 1;
	32909 : 1;
	32910 : 1;
	32911 : 1;
	32912 : 1;
	32913 : 1;
	32914 : 1;
	32915 : 1;
	32916 : 1;
	32917 : 1;
	32918 : 1;
	32919 : 1;
	32920 : 1;
	32921 : 1;
	32922 : 0;
	32923 : 0;
	32924 : 0;
	32925 : 1;
	32926 : 0;
	32927 : 1;
	32928 : 1;
	32929 : 1;
	32930 : 1;
	32931 : 0;
	32932 : 0;
	32933 : 0;
	32934 : 0;
	32935 : 1;
	32936 : 0;
	32937 : 1;
	32938 : 1;
	32939 : 1;
	32940 : 1;
	32941 : 1;
	32942 : 0;
	32943 : 0;
	32944 : 0;
	32945 : 0;
	32946 : 0;
	32947 : 1;
	32948 : 0;
	32949 : 0;
	32950 : 0;
	32951 : 1;
	32952 : 0;
	32953 : 1;
	32954 : 1;
	32955 : 0;
	32956 : 0;
	32957 : 0;
	32958 : 1;
	32959 : 1;
	32960 : 1;
	32961 : 0;
	32962 : 0;
	32963 : 0;
	32964 : 0;
	32965 : 1;
	32966 : 1;
	32967 : 0;
	32968 : 0;
	32969 : 0;
	32970 : 0;
	32971 : 0;
	32972 : 0;
	32973 : 0;
	32974 : 0;
	32975 : 0;
	32976 : 1;
	32977 : 0;
	32978 : 1;
	32979 : 0;
	32980 : 1;
	32981 : 0;
	32982 : 1;
	32983 : 0;
	32984 : 1;
	32985 : 1;
	32986 : 0;
	32987 : 0;
	32988 : 0;
	32989 : 0;
	32990 : 1;
	32991 : 0;
	32992 : 1;
	32993 : 1;
	32994 : 1;
	32995 : 1;
	32996 : 0;
	32997 : 0;
	32998 : 1;
	32999 : 1;
	33000 : 1;
	33001 : 1;
	33002 : 1;
	33003 : 1;
	33004 : 1;
	33005 : 1;
	33006 : 1;
	33007 : 1;
	33008 : 1;
	33009 : 0;
	33010 : 1;
	33011 : 1;
	33012 : 1;
	33013 : 0;
	33014 : 1;
	33015 : 0;
	33016 : 1;
	33017 : 1;
	33018 : 1;
	33019 : 1;
	33020 : 1;
	33021 : 0;
	33022 : 0;
	33023 : 0;
	33024 : 0;
	33025 : 1;
	33026 : 1;
	33027 : 0;
	33028 : 0;
	33029 : 0;
	33030 : 0;
	33031 : 0;
	33032 : 1;
	33033 : 1;
	33034 : 1;
	33035 : 1;
	33036 : 0;
	33037 : 0;
	33038 : 1;
	33039 : 0;
	33040 : 1;
	33041 : 0;
	33042 : 1;
	33043 : 1;
	33044 : 0;
	33045 : 0;
	33046 : 1;
	33047 : 0;
	33048 : 0;
	33049 : 0;
	33050 : 0;
	33051 : 0;
	33052 : 1;
	33053 : 1;
	33054 : 1;
	33055 : 0;
	33056 : 0;
	33057 : 0;
	33058 : 0;
	33059 : 0;
	33060 : 1;
	33061 : 0;
	33062 : 1;
	33063 : 0;
	33064 : 1;
	33065 : 0;
	33066 : 1;
	33067 : 0;
	33068 : 1;
	33069 : 1;
	33070 : 0;
	33071 : 1;
	33072 : 1;
	33073 : 0;
	33074 : 0;
	33075 : 0;
	33076 : 0;
	33077 : 0;
	33078 : 1;
	33079 : 1;
	33080 : 1;
	33081 : 1;
	33082 : 1;
	33083 : 1;
	33084 : 1;
	33085 : 1;
	33086 : 1;
	33087 : 1;
	33088 : 1;
	33089 : 1;
	33090 : 1;
	33091 : 1;
	33092 : 1;
	33093 : 1;
	33094 : 1;
	33095 : 1;
	33096 : 1;
	33097 : 1;
	33098 : 1;
	33099 : 1;
	33100 : 1;
	33101 : 1;
	33102 : 1;
	33103 : 1;
	33104 : 1;
	33105 : 1;
	33106 : 1;
	33107 : 1;
	33108 : 1;
	33109 : 1;
	33110 : 1;
	33111 : 1;
	33112 : 1;
	33113 : 1;
	33114 : 1;
	33115 : 1;
	33116 : 1;
	33117 : 1;
	33118 : 1;
	33119 : 1;
	33120 : 1;
	33121 : 1;
	33122 : 1;
	33123 : 1;
	33124 : 1;
	33125 : 1;
	33126 : 1;
	33127 : 1;
	33128 : 1;
	33129 : 1;
	33130 : 1;
	33131 : 1;
	33132 : 1;
	33133 : 1;
	33134 : 1;
	33135 : 1;
	33136 : 1;
	33137 : 1;
	33138 : 1;
	33139 : 1;
	33140 : 1;
	33141 : 1;
	33142 : 1;
	33143 : 1;
	33144 : 1;
	33145 : 1;
	33146 : 1;
	33147 : 1;
	33148 : 1;
	33149 : 1;
	33150 : 1;
	33151 : 1;
	33152 : 1;
	33153 : 1;
	33154 : 1;
	33155 : 1;
	33156 : 1;
	33157 : 1;
	33158 : 1;
	33159 : 1;
	33160 : 1;
	33161 : 1;
	33162 : 1;
	33163 : 1;
	33164 : 1;
	33165 : 1;
	33166 : 1;
	33167 : 1;
	33168 : 1;
	33169 : 1;
	33170 : 1;
	33171 : 1;
	33172 : 1;
	33173 : 1;
	33174 : 0;
	33175 : 1;
	33176 : 1;
	33177 : 1;
	33178 : 1;
	33179 : 1;
	33180 : 1;
	33181 : 1;
	33182 : 1;
	33183 : 1;
	33184 : 1;
	33185 : 1;
	33186 : 1;
	33187 : 1;
	33188 : 1;
	33189 : 1;
	33190 : 1;
	33191 : 1;
	33192 : 1;
	33193 : 1;
	33194 : 1;
	33195 : 1;
	33196 : 1;
	33197 : 1;
	33198 : 1;
	33199 : 1;
	33200 : 1;
	33201 : 1;
	33202 : 1;
	33203 : 1;
	33204 : 1;
	33205 : 1;
	33206 : 1;
	33207 : 1;
	33208 : 1;
	33209 : 1;
	33210 : 1;
	33211 : 1;
	33212 : 1;
	33213 : 1;
	33214 : 1;
	33215 : 1;
	33216 : 1;
	33217 : 1;
	33218 : 1;
	33219 : 1;
	33220 : 1;
	33221 : 1;
	33222 : 1;
	33223 : 1;
	33224 : 1;
	33225 : 1;
	33226 : 1;
	33227 : 1;
	33228 : 1;
	33229 : 1;
	33230 : 1;
	33231 : 1;
	33232 : 1;
	33233 : 1;
	33234 : 1;
	33235 : 1;
	33236 : 1;
	33237 : 1;
	33238 : 1;
	33239 : 1;
	33240 : 1;
	33241 : 1;
	33242 : 1;
	33243 : 1;
	33244 : 1;
	33245 : 1;
	33246 : 1;
	33247 : 1;
	33248 : 1;
	33249 : 1;
	33250 : 1;
	33251 : 1;
	33252 : 1;
	33253 : 1;
	33254 : 1;
	33255 : 1;
	33256 : 1;
	33257 : 1;
	33258 : 1;
	33259 : 1;
	33260 : 1;
	33261 : 1;
	33262 : 1;
	33263 : 1;
	33264 : 1;
	33265 : 1;
	33266 : 1;
	33267 : 1;
	33268 : 1;
	33269 : 1;
	33270 : 1;
	33271 : 0;
	33272 : 1;
	33273 : 1;
	33274 : 1;
	33275 : 1;
	33276 : 1;
	33277 : 1;
	33278 : 1;
	33279 : 1;
	33280 : 1;
	33281 : 1;
	33282 : 1;
	33283 : 1;
	33284 : 1;
	33285 : 1;
	33286 : 1;
	33287 : 1;
	33288 : 1;
	33289 : 1;
	33290 : 1;
	33291 : 1;
	33292 : 1;
	33293 : 1;
	33294 : 1;
	33295 : 1;
	33296 : 1;
	33297 : 1;
	33298 : 1;
	33299 : 1;
	33300 : 1;
	33301 : 1;
	33302 : 1;
	33303 : 1;
	33304 : 1;
	33305 : 1;
	33306 : 1;
	33307 : 1;
	33308 : 1;
	33309 : 1;
	33310 : 1;
	33311 : 1;
	33312 : 1;
	33313 : 1;
	33314 : 1;
	33315 : 1;
	33316 : 1;
	33317 : 0;
	33318 : 1;
	33319 : 1;
	33320 : 1;
	33321 : 1;
	33322 : 1;
	33323 : 1;
	33324 : 1;
	33325 : 1;
	33326 : 1;
	33327 : 1;
	33328 : 1;
	33329 : 1;
	33330 : 1;
	33331 : 1;
	33332 : 1;
	33333 : 1;
	33334 : 1;
	33335 : 1;
	33336 : 1;
	33337 : 1;
	33338 : 1;
	33339 : 1;
	33340 : 1;
	33341 : 1;
	33342 : 1;
	33343 : 1;
	33344 : 1;
	33345 : 1;
	33346 : 1;
	33347 : 1;
	33348 : 1;
	33349 : 1;
	33350 : 1;
	33351 : 1;
	33352 : 1;
	33353 : 1;
	33354 : 1;
	33355 : 1;
	33356 : 1;
	33357 : 1;
	33358 : 1;
	33359 : 1;
	33360 : 1;
	33361 : 1;
	33362 : 1;
	33363 : 1;
	33364 : 1;
	33365 : 1;
	33366 : 1;
	33367 : 1;
	33368 : 1;
	33369 : 1;
	33370 : 1;
	33371 : 1;
	33372 : 1;
	33373 : 1;
	33374 : 1;
	33375 : 1;
	33376 : 1;
	33377 : 1;
	33378 : 1;
	33379 : 1;
	33380 : 1;
	33381 : 1;
	33382 : 1;
	33383 : 1;
	33384 : 1;
	33385 : 1;
	33386 : 1;
	33387 : 1;
	33388 : 1;
	33389 : 1;
	33390 : 1;
	33391 : 1;
	33392 : 1;
	33393 : 1;
	33394 : 1;
	33395 : 1;
	33396 : 1;
	33397 : 1;
	33398 : 1;
	33399 : 1;
	33400 : 1;
	33401 : 1;
	33402 : 1;
	33403 : 1;
	33404 : 1;
	33405 : 1;
	33406 : 1;
	33407 : 1;
	33408 : 1;
	33409 : 1;
	33410 : 1;
	33411 : 0;
	33412 : 0;
	33413 : 0;
	33414 : 1;
	33415 : 1;
	33416 : 1;
	33417 : 1;
	33418 : 1;
	33419 : 1;
	33420 : 1;
	33421 : 1;
	33422 : 1;
	33423 : 1;
	33424 : 1;
	33425 : 1;
	33426 : 1;
	33427 : 1;
	33428 : 1;
	33429 : 1;
	33430 : 1;
	33431 : 1;
	33432 : 1;
	33433 : 1;
	33434 : 1;
	33435 : 1;
	33436 : 1;
	33437 : 1;
	33438 : 1;
	33439 : 1;
	33440 : 1;
	33441 : 1;
	33442 : 1;
	33443 : 1;
	33444 : 1;
	33445 : 1;
	33446 : 1;
	33447 : 1;
	33448 : 1;
	33449 : 1;
	33450 : 1;
	33451 : 1;
	33452 : 1;
	33453 : 1;
	33454 : 1;
	33455 : 1;
	33456 : 1;
	33457 : 1;
	33458 : 1;
	33459 : 1;
	33460 : 1;
	33461 : 1;
	33462 : 1;
	33463 : 1;
	33464 : 1;
	33465 : 1;
	33466 : 1;
	33467 : 1;
	33468 : 1;
	33469 : 1;
	33470 : 1;
	33471 : 1;
	33472 : 1;
	33473 : 1;
	33474 : 1;
	33475 : 1;
	33476 : 1;
	33477 : 1;
	33478 : 1;
	33479 : 1;
	33480 : 1;
	33481 : 1;
	33482 : 1;
	33483 : 1;
	33484 : 1;
	33485 : 1;
	33486 : 1;
	33487 : 1;
	33488 : 1;
	33489 : 1;
	33490 : 1;
	33491 : 1;
	33492 : 1;
	33493 : 1;
	33494 : 1;
	33495 : 1;
	33496 : 1;
	33497 : 1;
	33498 : 1;
	33499 : 1;
	33500 : 1;
	33501 : 1;
	33502 : 1;
	33503 : 1;
	33504 : 1;
	33505 : 1;
	33506 : 0;
	33507 : 0;
	33508 : 0;
	33509 : 0;
	33510 : 0;
	33511 : 1;
	33512 : 1;
	33513 : 1;
	33514 : 1;
	33515 : 1;
	33516 : 1;
	33517 : 1;
	33518 : 1;
	33519 : 1;
	33520 : 1;
	33521 : 1;
	33522 : 1;
	33523 : 1;
	33524 : 1;
	33525 : 1;
	33526 : 1;
	33527 : 1;
	33528 : 1;
	33529 : 1;
	33530 : 1;
	33531 : 1;
	33532 : 1;
	33533 : 1;
	33534 : 1;
	33535 : 1;
	33536 : 1;
	33537 : 1;
	33538 : 1;
	33539 : 1;
	33540 : 1;
	33541 : 1;
	33542 : 1;
	33543 : 1;
	33544 : 1;
	33545 : 1;
	33546 : 1;
	33547 : 1;
	33548 : 1;
	33549 : 1;
	33550 : 1;
	33551 : 1;
	33552 : 0;
	33553 : 0;
	33554 : 0;
	33555 : 0;
	33556 : 0;
	33557 : 1;
	33558 : 1;
	33559 : 1;
	33560 : 1;
	33561 : 1;
	33562 : 1;
	33563 : 1;
	33564 : 1;
	33565 : 1;
	33566 : 1;
	33567 : 1;
	33568 : 1;
	33569 : 1;
	33570 : 1;
	33571 : 1;
	33572 : 1;
	33573 : 1;
	33574 : 1;
	33575 : 1;
	33576 : 1;
	33577 : 1;
	33578 : 1;
	33579 : 1;
	33580 : 1;
	33581 : 1;
	33582 : 1;
	33583 : 1;
	33584 : 1;
	33585 : 1;
	33586 : 1;
	33587 : 1;
	33588 : 1;
	33589 : 1;
	33590 : 1;
	33591 : 1;
	33592 : 1;
	33593 : 1;
	33594 : 1;
	33595 : 1;
	33596 : 1;
	33597 : 1;
	33598 : 1;
	33599 : 1;
	33600 : 1;
	33601 : 1;
	33602 : 1;
	33603 : 1;
	33604 : 1;
	33605 : 1;
	33606 : 1;
	33607 : 1;
	33608 : 1;
	33609 : 1;
	33610 : 1;
	33611 : 1;
	33612 : 1;
	33613 : 1;
	33614 : 1;
	33615 : 1;
	33616 : 1;
	33617 : 1;
	33618 : 1;
	33619 : 1;
	33620 : 1;
	33621 : 1;
	33622 : 1;
	33623 : 1;
	33624 : 1;
	33625 : 1;
	33626 : 1;
	33627 : 1;
	33628 : 1;
	33629 : 1;
	33630 : 1;
	33631 : 1;
	33632 : 1;
	33633 : 1;
	33634 : 1;
	33635 : 1;
	33636 : 1;
	33637 : 1;
	33638 : 1;
	33639 : 1;
	33640 : 1;
	33641 : 1;
	33642 : 1;
	33643 : 1;
	33644 : 1;
	33645 : 1;
	33646 : 1;
	33647 : 1;
	33648 : 1;
	33649 : 1;
	33650 : 1;
	33651 : 1;
	33652 : 1;
	33653 : 1;
	33654 : 1;
	33655 : 1;
	33656 : 1;
	33657 : 1;
	33658 : 1;
	33659 : 1;
	33660 : 1;
	33661 : 1;
	33662 : 1;
	33663 : 1;
	33664 : 1;
	33665 : 1;
	33666 : 1;
	33667 : 1;
	33668 : 1;
	33669 : 1;
	33670 : 1;
	33671 : 1;
	33672 : 1;
	33673 : 1;
	33674 : 1;
	33675 : 1;
	33676 : 1;
	33677 : 1;
	33678 : 1;
	33679 : 1;
	33680 : 1;
	33681 : 1;
	33682 : 1;
	33683 : 1;
	33684 : 1;
	33685 : 1;
	33686 : 1;
	33687 : 1;
	33688 : 1;
	33689 : 1;
	33690 : 1;
	33691 : 1;
	33692 : 1;
	33693 : 1;
	33694 : 1;
	33695 : 1;
	33696 : 1;
	33697 : 1;
	33698 : 1;
	33699 : 1;
	33700 : 1;
	33701 : 1;
	33702 : 1;
	33703 : 1;
	33704 : 1;
	33705 : 1;
	33706 : 1;
	33707 : 1;
	33708 : 1;
	33709 : 1;
	33710 : 1;
	33711 : 1;
	33712 : 1;
	33713 : 1;
	33714 : 1;
	33715 : 1;
	33716 : 1;
	33717 : 1;
	33718 : 1;
	33719 : 1;
	33720 : 1;
	33721 : 1;
	33722 : 1;
	33723 : 1;
	33724 : 1;
	33725 : 1;
	33726 : 1;
	33727 : 1;
	33728 : 1;
	33729 : 1;
	33730 : 1;
	33731 : 1;
	33732 : 1;
	33733 : 1;
	33734 : 1;
	33735 : 1;
	33736 : 1;
	33737 : 1;
	33738 : 1;
	33739 : 1;
	33740 : 1;
	33741 : 1;
	33742 : 1;
	33743 : 1;
	33744 : 1;
	33745 : 1;
	33746 : 1;
	33747 : 1;
	33748 : 1;
	33749 : 1;
	33750 : 1;
	33751 : 1;
	33752 : 1;
	33753 : 1;
	33754 : 1;
	33755 : 1;
	33756 : 1;
	33757 : 1;
	33758 : 1;
	33759 : 1;
	33760 : 1;
	33761 : 1;
	33762 : 1;
	33763 : 1;
	33764 : 1;
	33765 : 1;
	33766 : 1;
	33767 : 1;
	33768 : 1;
	33769 : 1;
	33770 : 1;
	33771 : 1;
	33772 : 1;
	33773 : 1;
	33774 : 1;
	33775 : 1;
	33776 : 1;
	33777 : 1;
	33778 : 1;
	33779 : 1;
	33780 : 1;
	33781 : 1;
	33782 : 1;
	33783 : 1;
	33784 : 1;
	33785 : 1;
	33786 : 1;
	33787 : 1;
	33788 : 1;
	33789 : 1;
	33790 : 1;
	33791 : 1;
	33792 : 1;
	33793 : 1;
	33794 : 1;
	33795 : 1;
	33796 : 1;
	33797 : 1;
	33798 : 1;
	33799 : 1;
	33800 : 1;
	33801 : 1;
	33802 : 1;
	33803 : 1;
	33804 : 1;
	33805 : 1;
	33806 : 1;
	33807 : 1;
	33808 : 1;
	33809 : 1;
	33810 : 1;
	33811 : 1;
	33812 : 1;
	33813 : 1;
	33814 : 1;
	33815 : 1;
	33816 : 1;
	33817 : 1;
	33818 : 1;
	33819 : 1;
	33820 : 1;
	33821 : 1;
	33822 : 1;
	33823 : 1;
	33824 : 1;
	33825 : 1;
	33826 : 1;
	33827 : 1;
	33828 : 1;
	33829 : 1;
	33830 : 1;
	33831 : 1;
	33832 : 1;
	33833 : 1;
	33834 : 1;
	33835 : 1;
	33836 : 1;
	33837 : 1;
	33838 : 1;
	33839 : 1;
	33840 : 1;
	33841 : 1;
	33842 : 1;
	33843 : 1;
	33844 : 1;
	33845 : 1;
	33846 : 1;
	33847 : 1;
	33848 : 1;
	33849 : 1;
	33850 : 1;
	33851 : 1;
	33852 : 1;
	33853 : 1;
	33854 : 1;
	33855 : 1;
	33856 : 1;
	33857 : 1;
	33858 : 1;
	33859 : 1;
	33860 : 1;
	33861 : 1;
	33862 : 1;
	33863 : 1;
	33864 : 1;
	33865 : 1;
	33866 : 1;
	33867 : 1;
	33868 : 1;
	33869 : 1;
	33870 : 1;
	33871 : 1;
	33872 : 1;
	33873 : 1;
	33874 : 1;
	33875 : 1;
	33876 : 1;
	33877 : 1;
	33878 : 1;
	33879 : 1;
	33880 : 1;
	33881 : 1;
	33882 : 1;
	33883 : 1;
	33884 : 1;
	33885 : 1;
	33886 : 1;
	33887 : 1;
	33888 : 1;
	33889 : 1;
	33890 : 1;
	33891 : 1;
	33892 : 1;
	33893 : 1;
	33894 : 1;
	33895 : 1;
	33896 : 1;
	33897 : 1;
	33898 : 1;
	33899 : 1;
	33900 : 1;
	33901 : 1;
	33902 : 1;
	33903 : 1;
	33904 : 1;
	33905 : 1;
	33906 : 1;
	33907 : 1;
	33908 : 1;
	33909 : 1;
	33910 : 1;
	33911 : 1;
	33912 : 1;
	33913 : 1;
	33914 : 1;
	33915 : 1;
	33916 : 1;
	33917 : 1;
	33918 : 1;
	33919 : 1;
	33920 : 1;
	33921 : 1;
	33922 : 1;
	33923 : 1;
	33924 : 1;
	33925 : 1;
	33926 : 1;
	33927 : 1;
	33928 : 1;
	33929 : 1;
	33930 : 1;
	33931 : 1;
	33932 : 1;
	33933 : 1;
	33934 : 1;
	33935 : 1;
	33936 : 1;
	33937 : 1;
	33938 : 1;
	33939 : 1;
	33940 : 1;
	33941 : 1;
	33942 : 1;
	33943 : 1;
	33944 : 1;
	33945 : 1;
	33946 : 1;
	33947 : 1;
	33948 : 1;
	33949 : 1;
	33950 : 1;
	33951 : 1;
	33952 : 1;
	33953 : 1;
	33954 : 1;
	33955 : 1;
	33956 : 1;
	33957 : 1;
	33958 : 1;
	33959 : 1;
	33960 : 1;
	33961 : 1;
	33962 : 1;
	33963 : 1;
	33964 : 1;
	33965 : 1;
	33966 : 1;
	33967 : 1;
	33968 : 1;
	33969 : 1;
	33970 : 1;
	33971 : 1;
	33972 : 1;
	33973 : 1;
	33974 : 1;
	33975 : 1;
	33976 : 1;
	33977 : 1;
	33978 : 1;
	33979 : 1;
	33980 : 1;
	33981 : 1;
	33982 : 1;
	33983 : 1;
	33984 : 1;
	33985 : 1;
	33986 : 1;
	33987 : 1;
	33988 : 1;
	33989 : 1;
	33990 : 1;
	33991 : 1;
	33992 : 1;
	33993 : 1;
	33994 : 1;
	33995 : 1;
	33996 : 1;
	33997 : 1;
	33998 : 1;
	33999 : 1;
	34000 : 1;
	34001 : 1;
	34002 : 1;
	34003 : 1;
	34004 : 1;
	34005 : 1;
	34006 : 1;
	34007 : 1;
	34008 : 1;
	34009 : 1;
	34010 : 1;
	34011 : 1;
	34012 : 1;
	34013 : 1;
	34014 : 1;
	34015 : 1;
	34016 : 1;
	34017 : 1;
	34018 : 1;
	34019 : 1;
	34020 : 1;
	34021 : 1;
	34022 : 1;
	34023 : 1;
	34024 : 1;
	34025 : 1;
	34026 : 1;
	34027 : 1;
	34028 : 1;
	34029 : 1;
	34030 : 1;
	34031 : 1;
	34032 : 1;
	34033 : 1;
	34034 : 1;
	34035 : 1;
	34036 : 1;
	34037 : 1;
	34038 : 1;
	34039 : 1;
	34040 : 1;
	34041 : 1;
	34042 : 1;
	34043 : 1;
	34044 : 1;
	34045 : 1;
	34046 : 1;
	34047 : 1;
	34048 : 1;
	34049 : 1;
	34050 : 1;
	34051 : 1;
	34052 : 1;
	34053 : 1;
	34054 : 1;
	34055 : 1;
	34056 : 1;
	34057 : 1;
	34058 : 1;
	34059 : 1;
	34060 : 1;
	34061 : 1;
	34062 : 1;
	34063 : 1;
	34064 : 1;
	34065 : 1;
	34066 : 1;
	34067 : 1;
	34068 : 1;
	34069 : 1;
	34070 : 1;
	34071 : 1;
	34072 : 1;
	34073 : 1;
	34074 : 1;
	34075 : 1;
	34076 : 1;
	34077 : 1;
	34078 : 1;
	34079 : 1;
	34080 : 1;
	34081 : 1;
	34082 : 1;
	34083 : 1;
	34084 : 1;
	34085 : 1;
	34086 : 1;
	34087 : 1;
	34088 : 1;
	34089 : 1;
	34090 : 1;
	34091 : 1;
	34092 : 1;
	34093 : 1;
	34094 : 1;
	34095 : 1;
	34096 : 1;
	34097 : 1;
	34098 : 1;
	34099 : 1;
	34100 : 1;
	34101 : 1;
	34102 : 1;
	34103 : 1;
	34104 : 1;
	34105 : 1;
	34106 : 1;
	34107 : 1;
	34108 : 1;
	34109 : 1;
	34110 : 1;
	34111 : 1;
	34112 : 1;
	34113 : 1;
	34114 : 1;
	34115 : 1;
	34116 : 1;
	34117 : 1;
	34118 : 1;
	34119 : 1;
	34120 : 1;
	34121 : 1;
	34122 : 1;
	34123 : 1;
	34124 : 1;
	34125 : 1;
	34126 : 1;
	34127 : 1;
	34128 : 1;
	34129 : 1;
	34130 : 1;
	34131 : 1;
	34132 : 1;
	34133 : 1;
	34134 : 1;
	34135 : 1;
	34136 : 1;
	34137 : 1;
	34138 : 1;
	34139 : 1;
	34140 : 1;
	34141 : 1;
	34142 : 1;
	34143 : 1;
	34144 : 1;
	34145 : 1;
	34146 : 1;
	34147 : 1;
	34148 : 1;
	34149 : 1;
	34150 : 1;
	34151 : 1;
	34152 : 1;
	34153 : 1;
	34154 : 1;
	34155 : 1;
	34156 : 1;
	34157 : 1;
	34158 : 1;
	34159 : 1;
	34160 : 1;
	34161 : 1;
	34162 : 1;
	34163 : 1;
	34164 : 1;
	34165 : 1;
	34166 : 1;
	34167 : 1;
	34168 : 1;
	34169 : 1;
	34170 : 1;
	34171 : 1;
	34172 : 1;
	34173 : 1;
	34174 : 1;
	34175 : 1;
	34176 : 1;
	34177 : 1;
	34178 : 1;
	34179 : 1;
	34180 : 1;
	34181 : 1;
	34182 : 1;
	34183 : 1;
	34184 : 1;
	34185 : 1;
	34186 : 1;
	34187 : 1;
	34188 : 1;
	34189 : 1;
	34190 : 1;
	34191 : 1;
	34192 : 1;
	34193 : 1;
	34194 : 1;
	34195 : 1;
	34196 : 1;
	34197 : 1;
	34198 : 1;
	34199 : 1;
	34200 : 1;
	34201 : 1;
	34202 : 1;
	34203 : 1;
	34204 : 1;
	34205 : 1;
	34206 : 1;
	34207 : 1;
	34208 : 1;
	34209 : 1;
	34210 : 1;
	34211 : 1;
	34212 : 1;
	34213 : 1;
	34214 : 1;
	34215 : 1;
	34216 : 1;
	34217 : 1;
	34218 : 1;
	34219 : 1;
	34220 : 1;
	34221 : 1;
	34222 : 1;
	34223 : 1;
	34224 : 1;
	34225 : 1;
	34226 : 1;
	34227 : 1;
	34228 : 1;
	34229 : 1;
	34230 : 1;
	34231 : 1;
	34232 : 1;
	34233 : 1;
	34234 : 1;
	34235 : 1;
	34236 : 1;
	34237 : 1;
	34238 : 1;
	34239 : 1;
	34240 : 1;
	34241 : 1;
	34242 : 1;
	34243 : 1;
	34244 : 1;
	34245 : 1;
	34246 : 1;
	34247 : 1;
	34248 : 1;
	34249 : 1;
	34250 : 1;
	34251 : 1;
	34252 : 1;
	34253 : 1;
	34254 : 1;
	34255 : 1;
	34256 : 1;
	34257 : 1;
	34258 : 1;
	34259 : 1;
	34260 : 1;
	34261 : 1;
	34262 : 1;
	34263 : 1;
	34264 : 1;
	34265 : 1;
	34266 : 1;
	34267 : 1;
	34268 : 1;
	34269 : 1;
	34270 : 1;
	34271 : 1;
	34272 : 1;
	34273 : 1;
	34274 : 1;
	34275 : 1;
	34276 : 1;
	34277 : 1;
	34278 : 1;
	34279 : 1;
	34280 : 1;
	34281 : 1;
	34282 : 1;
	34283 : 1;
	34284 : 1;
	34285 : 1;
	34286 : 1;
	34287 : 1;
	34288 : 1;
	34289 : 1;
	34290 : 1;
	34291 : 1;
	34292 : 1;
	34293 : 1;
	34294 : 1;
	34295 : 1;
	34296 : 1;
	34297 : 1;
	34298 : 1;
	34299 : 1;
	34300 : 1;
	34301 : 1;
	34302 : 1;
	34303 : 1;
	34304 : 1;
	34305 : 1;
	34306 : 1;
	34307 : 1;
	34308 : 1;
	34309 : 1;
	34310 : 1;
	34311 : 1;
	34312 : 1;
	34313 : 1;
	34314 : 1;
	34315 : 1;
	34316 : 1;
	34317 : 1;
	34318 : 1;
	34319 : 1;
	34320 : 1;
	34321 : 1;
	34322 : 1;
	34323 : 1;
	34324 : 1;
	34325 : 1;
	34326 : 1;
	34327 : 1;
	34328 : 1;
	34329 : 1;
	34330 : 1;
	34331 : 1;
	34332 : 1;
	34333 : 1;
	34334 : 1;
	34335 : 1;
	34336 : 1;
	34337 : 1;
	34338 : 1;
	34339 : 1;
	34340 : 1;
	34341 : 1;
	34342 : 1;
	34343 : 1;
	34344 : 1;
	34345 : 1;
	34346 : 1;
	34347 : 1;
	34348 : 1;
	34349 : 1;
	34350 : 1;
	34351 : 1;
	34352 : 1;
	34353 : 1;
	34354 : 1;
	34355 : 1;
	34356 : 1;
	34357 : 1;
	34358 : 1;
	34359 : 1;
	34360 : 1;
	34361 : 1;
	34362 : 1;
	34363 : 1;
	34364 : 1;
	34365 : 1;
	34366 : 1;
	34367 : 1;
	34368 : 1;
	34369 : 1;
	34370 : 1;
	34371 : 1;
	34372 : 1;
	34373 : 1;
	34374 : 1;
	34375 : 1;
	34376 : 1;
	34377 : 1;
	34378 : 1;
	34379 : 1;
	34380 : 1;
	34381 : 1;
	34382 : 1;
	34383 : 1;
	34384 : 1;
	34385 : 1;
	34386 : 1;
	34387 : 1;
	34388 : 1;
	34389 : 1;
	34390 : 1;
	34391 : 1;
	34392 : 1;
	34393 : 1;
	34394 : 1;
	34395 : 1;
	34396 : 1;
	34397 : 1;
	34398 : 1;
	34399 : 1;
	34400 : 1;
	34401 : 1;
	34402 : 1;
	34403 : 1;
	34404 : 1;
	34405 : 1;
	34406 : 1;
	34407 : 1;
	34408 : 1;
	34409 : 1;
	34410 : 1;
	34411 : 1;
	34412 : 1;
	34413 : 1;
	34414 : 1;
	34415 : 1;
	34416 : 1;
	34417 : 1;
	34418 : 1;
	34419 : 1;
	34420 : 1;
	34421 : 1;
	34422 : 1;
	34423 : 1;
	34424 : 1;
	34425 : 1;
	34426 : 1;
	34427 : 1;
	34428 : 1;
	34429 : 1;
	34430 : 1;
	34431 : 1;
	34432 : 1;
	34433 : 1;
	34434 : 1;
	34435 : 1;
	34436 : 1;
	34437 : 1;
	34438 : 1;
	34439 : 1;
	34440 : 1;
	34441 : 1;
	34442 : 1;
	34443 : 1;
	34444 : 1;
	34445 : 1;
	34446 : 1;
	34447 : 1;
	34448 : 1;
	34449 : 1;
	34450 : 1;
	34451 : 1;
	34452 : 1;
	34453 : 1;
	34454 : 1;
	34455 : 1;
	34456 : 1;
	34457 : 1;
	34458 : 1;
	34459 : 1;
	34460 : 1;
	34461 : 1;
	34462 : 1;
	34463 : 1;
	34464 : 1;
	34465 : 1;
	34466 : 1;
	34467 : 1;
	34468 : 1;
	34469 : 1;
	34470 : 1;
	34471 : 1;
	34472 : 1;
	34473 : 1;
	34474 : 1;
	34475 : 1;
	34476 : 1;
	34477 : 1;
	34478 : 1;
	34479 : 1;
	34480 : 1;
	34481 : 1;
	34482 : 1;
	34483 : 1;
	34484 : 1;
	34485 : 1;
	34486 : 1;
	34487 : 1;
	34488 : 1;
	34489 : 1;
	34490 : 1;
	34491 : 1;
	34492 : 1;
	34493 : 1;
	34494 : 1;
	34495 : 1;
	34496 : 1;
	34497 : 1;
	34498 : 1;
	34499 : 1;
	34500 : 1;
	34501 : 1;
	34502 : 1;
	34503 : 1;
	34504 : 1;
	34505 : 1;
	34506 : 1;
	34507 : 1;
	34508 : 1;
	34509 : 1;
	34510 : 1;
	34511 : 1;
	34512 : 1;
	34513 : 1;
	34514 : 1;
	34515 : 1;
	34516 : 1;
	34517 : 1;
	34518 : 1;
	34519 : 1;
	34520 : 1;
	34521 : 1;
	34522 : 1;
	34523 : 1;
	34524 : 1;
	34525 : 1;
	34526 : 1;
	34527 : 1;
	34528 : 1;
	34529 : 1;
	34530 : 1;
	34531 : 1;
	34532 : 1;
	34533 : 1;
	34534 : 1;
	34535 : 1;
	34536 : 1;
	34537 : 1;
	34538 : 1;
	34539 : 1;
	34540 : 1;
	34541 : 1;
	34542 : 1;
	34543 : 1;
	34544 : 1;
	34545 : 1;
	34546 : 1;
	34547 : 1;
	34548 : 1;
	34549 : 1;
	34550 : 1;
	34551 : 1;
	34552 : 1;
	34553 : 1;
	34554 : 1;
	34555 : 1;
	34556 : 1;
	34557 : 1;
	34558 : 1;
	34559 : 1;
	34560 : 1;
	34561 : 1;
	34562 : 1;
	34563 : 1;
	34564 : 1;
	34565 : 1;
	34566 : 1;
	34567 : 1;
	34568 : 1;
	34569 : 1;
	34570 : 1;
	34571 : 1;
	34572 : 1;
	34573 : 1;
	34574 : 1;
	34575 : 1;
	34576 : 1;
	34577 : 1;
	34578 : 1;
	34579 : 1;
	34580 : 1;
	34581 : 1;
	34582 : 1;
	34583 : 1;
	34584 : 1;
	34585 : 1;
	34586 : 1;
	34587 : 1;
	34588 : 1;
	34589 : 1;
	34590 : 1;
	34591 : 1;
	34592 : 1;
	34593 : 1;
	34594 : 1;
	34595 : 1;
	34596 : 1;
	34597 : 1;
	34598 : 1;
	34599 : 1;
	34600 : 1;
	34601 : 1;
	34602 : 1;
	34603 : 1;
	34604 : 1;
	34605 : 1;
	34606 : 1;
	34607 : 1;
	34608 : 1;
	34609 : 1;
	34610 : 1;
	34611 : 1;
	34612 : 1;
	34613 : 1;
	34614 : 1;
	34615 : 1;
	34616 : 1;
	34617 : 1;
	34618 : 1;
	34619 : 1;
	34620 : 1;
	34621 : 1;
	34622 : 1;
	34623 : 1;
	34624 : 1;
	34625 : 1;
	34626 : 1;
	34627 : 1;
	34628 : 1;
	34629 : 1;
	34630 : 1;
	34631 : 1;
	34632 : 1;
	34633 : 1;
	34634 : 1;
	34635 : 1;
	34636 : 1;
	34637 : 1;
	34638 : 1;
	34639 : 1;
	34640 : 1;
	34641 : 1;
	34642 : 1;
	34643 : 1;
	34644 : 1;
	34645 : 1;
	34646 : 1;
	34647 : 1;
	34648 : 1;
	34649 : 1;
	34650 : 1;
	34651 : 1;
	34652 : 1;
	34653 : 1;
	34654 : 1;
	34655 : 1;
	34656 : 1;
	34657 : 1;
	34658 : 1;
	34659 : 1;
	34660 : 1;
	34661 : 1;
	34662 : 1;
	34663 : 1;
	34664 : 1;
	34665 : 1;
	34666 : 1;
	34667 : 1;
	34668 : 1;
	34669 : 1;
	34670 : 1;
	34671 : 1;
	34672 : 1;
	34673 : 1;
	34674 : 1;
	34675 : 1;
	34676 : 1;
	34677 : 1;
	34678 : 1;
	34679 : 1;
	34680 : 1;
	34681 : 1;
	34682 : 1;
	34683 : 1;
	34684 : 1;
	34685 : 1;
	34686 : 1;
	34687 : 1;
	34688 : 1;
	34689 : 1;
	34690 : 1;
	34691 : 1;
	34692 : 1;
	34693 : 1;
	34694 : 1;
	34695 : 1;
	34696 : 1;
	34697 : 1;
	34698 : 1;
	34699 : 1;
	34700 : 1;
	34701 : 1;
	34702 : 1;
	34703 : 1;
	34704 : 1;
	34705 : 1;
	34706 : 1;
	34707 : 1;
	34708 : 1;
	34709 : 1;
	34710 : 1;
	34711 : 1;
	34712 : 1;
	34713 : 1;
	34714 : 1;
	34715 : 1;
	34716 : 1;
	34717 : 1;
	34718 : 1;
	34719 : 1;
	34720 : 1;
	34721 : 1;
	34722 : 1;
	34723 : 1;
	34724 : 1;
	34725 : 1;
	34726 : 1;
	34727 : 1;
	34728 : 1;
	34729 : 1;
	34730 : 1;
	34731 : 1;
	34732 : 1;
	34733 : 1;
	34734 : 1;
	34735 : 1;
	34736 : 1;
	34737 : 1;
	34738 : 1;
	34739 : 1;
	34740 : 1;
	34741 : 1;
	34742 : 1;
	34743 : 1;
	34744 : 1;
	34745 : 1;
	34746 : 1;
	34747 : 1;
	34748 : 1;
	34749 : 1;
	34750 : 1;
	34751 : 1;
	34752 : 1;
	34753 : 1;
	34754 : 1;
	34755 : 1;
	34756 : 1;
	34757 : 1;
	34758 : 1;
	34759 : 1;
	34760 : 1;
	34761 : 1;
	34762 : 1;
	34763 : 1;
	34764 : 1;
	34765 : 1;
	34766 : 1;
	34767 : 1;
	34768 : 1;
	34769 : 1;
	34770 : 1;
	34771 : 1;
	34772 : 1;
	34773 : 1;
	34774 : 1;
	34775 : 1;
	34776 : 1;
	34777 : 1;
	34778 : 1;
	34779 : 1;
	34780 : 1;
	34781 : 1;
	34782 : 1;
	34783 : 1;
	34784 : 1;
	34785 : 1;
	34786 : 1;
	34787 : 1;
	34788 : 1;
	34789 : 1;
	34790 : 1;
	34791 : 1;
	34792 : 1;
	34793 : 1;
	34794 : 1;
	34795 : 1;
	34796 : 1;
	34797 : 1;
	34798 : 1;
	34799 : 1;
	34800 : 1;
	34801 : 1;
	34802 : 1;
	34803 : 1;
	34804 : 1;
	34805 : 1;
	34806 : 1;
	34807 : 1;
	34808 : 1;
	34809 : 1;
	34810 : 1;
	34811 : 1;
	34812 : 1;
	34813 : 1;
	34814 : 1;
	34815 : 1;
	34816 : 1;
	34817 : 1;
	34818 : 1;
	34819 : 1;
	34820 : 1;
	34821 : 1;
	34822 : 1;
	34823 : 1;
	34824 : 1;
	34825 : 1;
	34826 : 1;
	34827 : 1;
	34828 : 1;
	34829 : 1;
	34830 : 1;
	34831 : 1;
	34832 : 1;
	34833 : 1;
	34834 : 1;
	34835 : 1;
	34836 : 1;
	34837 : 1;
	34838 : 1;
	34839 : 1;
	34840 : 1;
	34841 : 1;
	34842 : 1;
	34843 : 1;
	34844 : 1;
	34845 : 1;
	34846 : 1;
	34847 : 1;
	34848 : 1;
	34849 : 1;
	34850 : 1;
	34851 : 1;
	34852 : 1;
	34853 : 1;
	34854 : 1;
	34855 : 1;
	34856 : 1;
	34857 : 1;
	34858 : 1;
	34859 : 1;
	34860 : 1;
	34861 : 1;
	34862 : 1;
	34863 : 1;
	34864 : 1;
	34865 : 1;
	34866 : 1;
	34867 : 1;
	34868 : 1;
	34869 : 1;
	34870 : 1;
	34871 : 1;
	34872 : 1;
	34873 : 1;
	34874 : 1;
	34875 : 1;
	34876 : 1;
	34877 : 1;
	34878 : 1;
	34879 : 1;
	34880 : 1;
	34881 : 1;
	34882 : 1;
	34883 : 1;
	34884 : 1;
	34885 : 1;
	34886 : 1;
	34887 : 1;
	34888 : 1;
	34889 : 1;
	34890 : 1;
	34891 : 1;
	34892 : 1;
	34893 : 1;
	34894 : 1;
	34895 : 1;
	34896 : 1;
	34897 : 1;
	34898 : 1;
	34899 : 1;
	34900 : 1;
	34901 : 1;
	34902 : 1;
	34903 : 1;
	34904 : 1;
	34905 : 1;
	34906 : 1;
	34907 : 1;
	34908 : 1;
	34909 : 1;
	34910 : 1;
	34911 : 1;
	34912 : 1;
	34913 : 1;
	34914 : 1;
	34915 : 1;
	34916 : 1;
	34917 : 1;
	34918 : 1;
	34919 : 1;
	34920 : 1;
	34921 : 1;
	34922 : 1;
	34923 : 1;
	34924 : 1;
	34925 : 1;
	34926 : 1;
	34927 : 1;
	34928 : 1;
	34929 : 1;
	34930 : 1;
	34931 : 1;
	34932 : 1;
	34933 : 1;
	34934 : 1;
	34935 : 1;
	34936 : 1;
	34937 : 1;
	34938 : 1;
	34939 : 1;
	34940 : 1;
	34941 : 1;
	34942 : 1;
	34943 : 1;
	34944 : 1;
	34945 : 1;
	34946 : 1;
	34947 : 1;
	34948 : 1;
	34949 : 1;
	34950 : 1;
	34951 : 1;
	34952 : 1;
	34953 : 1;
	34954 : 1;
	34955 : 1;
	34956 : 1;
	34957 : 1;
	34958 : 1;
	34959 : 1;
	34960 : 1;
	34961 : 1;
	34962 : 1;
	34963 : 1;
	34964 : 1;
	34965 : 1;
	34966 : 1;
	34967 : 1;
	34968 : 1;
	34969 : 1;
	34970 : 1;
	34971 : 1;
	34972 : 1;
	34973 : 1;
	34974 : 1;
	34975 : 1;
	34976 : 1;
	34977 : 1;
	34978 : 1;
	34979 : 1;
	34980 : 1;
	34981 : 1;
	34982 : 1;
	34983 : 1;
	34984 : 1;
	34985 : 1;
	34986 : 1;
	34987 : 1;
	34988 : 1;
	34989 : 1;
	34990 : 1;
	34991 : 1;
	34992 : 1;
	34993 : 1;
	34994 : 1;
	34995 : 1;
	34996 : 1;
	34997 : 1;
	34998 : 1;
	34999 : 1;
	35000 : 1;
	35001 : 1;
	35002 : 1;
	35003 : 1;
	35004 : 1;
	35005 : 1;
	35006 : 1;
	35007 : 1;
	35008 : 1;
	35009 : 1;
	35010 : 1;
	35011 : 1;
	35012 : 1;
	35013 : 1;
	35014 : 1;
	35015 : 1;
	35016 : 1;
	35017 : 1;
	35018 : 1;
	35019 : 1;
	35020 : 1;
	35021 : 1;
	35022 : 1;
	35023 : 1;
	35024 : 1;
	35025 : 1;
	35026 : 1;
	35027 : 1;
	35028 : 1;
	35029 : 1;
	35030 : 1;
	35031 : 1;
	35032 : 1;
	35033 : 1;
	35034 : 1;
	35035 : 1;
	35036 : 1;
	35037 : 1;
	35038 : 1;
	35039 : 1;
	35040 : 1;
	35041 : 1;
	35042 : 1;
	35043 : 1;
	35044 : 1;
	35045 : 1;
	35046 : 1;
	35047 : 1;
	35048 : 1;
	35049 : 1;
	35050 : 1;
	35051 : 1;
	35052 : 1;
	35053 : 1;
	35054 : 1;
	35055 : 1;
	35056 : 1;
	35057 : 1;
	35058 : 1;
	35059 : 1;
	35060 : 1;
	35061 : 1;
	35062 : 1;
	35063 : 1;
	35064 : 1;
	35065 : 1;
	35066 : 1;
	35067 : 1;
	35068 : 1;
	35069 : 1;
	35070 : 1;
	35071 : 1;
	35072 : 1;
	35073 : 1;
	35074 : 1;
	35075 : 1;
	35076 : 1;
	35077 : 1;
	35078 : 1;
	35079 : 1;
	35080 : 1;
	35081 : 1;
	35082 : 1;
	35083 : 1;
	35084 : 1;
	35085 : 1;
	35086 : 1;
	35087 : 1;
	35088 : 1;
	35089 : 1;
	35090 : 1;
	35091 : 1;
	35092 : 1;
	35093 : 1;
	35094 : 1;
	35095 : 1;
	35096 : 1;
	35097 : 1;
	35098 : 1;
	35099 : 1;
	35100 : 1;
	35101 : 1;
	35102 : 1;
	35103 : 1;
	35104 : 1;
	35105 : 1;
	35106 : 1;
	35107 : 1;
	35108 : 1;
	35109 : 1;
	35110 : 1;
	35111 : 1;
	35112 : 1;
	35113 : 1;
	35114 : 1;
	35115 : 1;
	35116 : 1;
	35117 : 1;
	35118 : 1;
	35119 : 1;
	35120 : 1;
	35121 : 1;
	35122 : 1;
	35123 : 1;
	35124 : 1;
	35125 : 1;
	35126 : 1;
	35127 : 1;
	35128 : 1;
	35129 : 1;
	35130 : 1;
	35131 : 1;
	35132 : 1;
	35133 : 1;
	35134 : 1;
	35135 : 1;
	35136 : 1;
	35137 : 1;
	35138 : 1;
	35139 : 1;
	35140 : 1;
	35141 : 1;
	35142 : 1;
	35143 : 1;
	35144 : 1;
	35145 : 1;
	35146 : 1;
	35147 : 1;
	35148 : 1;
	35149 : 1;
	35150 : 1;
	35151 : 1;
	35152 : 1;
	35153 : 1;
	35154 : 1;
	35155 : 1;
	35156 : 1;
	35157 : 1;
	35158 : 1;
	35159 : 1;
	35160 : 1;
	35161 : 1;
	35162 : 1;
	35163 : 1;
	35164 : 1;
	35165 : 1;
	35166 : 1;
	35167 : 1;
	35168 : 1;
	35169 : 1;
	35170 : 1;
	35171 : 1;
	35172 : 1;
	35173 : 1;
	35174 : 1;
	35175 : 1;
	35176 : 1;
	35177 : 1;
	35178 : 1;
	35179 : 1;
	35180 : 1;
	35181 : 1;
	35182 : 1;
	35183 : 1;
	35184 : 1;
	35185 : 1;
	35186 : 1;
	35187 : 1;
	35188 : 1;
	35189 : 1;
	35190 : 1;
	35191 : 1;
	35192 : 1;
	35193 : 1;
	35194 : 1;
	35195 : 1;
	35196 : 1;
	35197 : 1;
	35198 : 1;
	35199 : 1;
	35200 : 1;
	35201 : 1;
	35202 : 1;
	35203 : 1;
	35204 : 1;
	35205 : 1;
	35206 : 1;
	35207 : 1;
	35208 : 1;
	35209 : 1;
	35210 : 1;
	35211 : 1;
	35212 : 1;
	35213 : 1;
	35214 : 1;
	35215 : 1;
	35216 : 1;
	35217 : 1;
	35218 : 1;
	35219 : 1;
	35220 : 1;
	35221 : 1;
	35222 : 1;
	35223 : 1;
	35224 : 1;
	35225 : 1;
	35226 : 1;
	35227 : 1;
	35228 : 1;
	35229 : 1;
	35230 : 1;
	35231 : 1;
	35232 : 1;
	35233 : 1;
	35234 : 1;
	35235 : 1;
	35236 : 1;
	35237 : 1;
	35238 : 1;
	35239 : 1;
	35240 : 1;
	35241 : 1;
	35242 : 1;
	35243 : 1;
	35244 : 1;
	35245 : 1;
	35246 : 1;
	35247 : 1;
	35248 : 1;
	35249 : 1;
	35250 : 1;
	35251 : 1;
	35252 : 1;
	35253 : 1;
	35254 : 1;
	35255 : 1;
	35256 : 1;
	35257 : 1;
	35258 : 1;
	35259 : 1;
	35260 : 1;
	35261 : 1;
	35262 : 1;
	35263 : 1;
	35264 : 1;
	35265 : 1;
	35266 : 1;
	35267 : 1;
	35268 : 1;
	35269 : 1;
	35270 : 1;
	35271 : 1;
	35272 : 1;
	35273 : 1;
	35274 : 1;
	35275 : 1;
	35276 : 1;
	35277 : 1;
	35278 : 1;
	35279 : 1;
	35280 : 1;
	35281 : 1;
	35282 : 1;
	35283 : 1;
	35284 : 1;
	35285 : 1;
	35286 : 1;
	35287 : 1;
	35288 : 1;
	35289 : 1;
	35290 : 1;
	35291 : 1;
	35292 : 1;
	35293 : 1;
	35294 : 1;
	35295 : 1;
	35296 : 1;
	35297 : 1;
	35298 : 1;
	35299 : 1;
	35300 : 1;
	35301 : 1;
	35302 : 1;
	35303 : 1;
	35304 : 1;
	35305 : 1;
	35306 : 1;
	35307 : 1;
	35308 : 1;
	35309 : 1;
	35310 : 1;
	35311 : 1;
	35312 : 1;
	35313 : 1;
	35314 : 1;
	35315 : 1;
	35316 : 1;
	35317 : 1;
	35318 : 1;
	35319 : 1;
	35320 : 1;
	35321 : 1;
	35322 : 1;
	35323 : 1;
	35324 : 1;
	35325 : 1;
	35326 : 1;
	35327 : 1;
	35328 : 1;
	35329 : 0;
	35330 : 0;
	35331 : 0;
	35332 : 1;
	35333 : 1;
	35334 : 0;
	35335 : 0;
	35336 : 0;
	35337 : 1;
	35338 : 1;
	35339 : 0;
	35340 : 1;
	35341 : 1;
	35342 : 1;
	35343 : 1;
	35344 : 1;
	35345 : 1;
	35346 : 1;
	35347 : 1;
	35348 : 1;
	35349 : 1;
	35350 : 1;
	35351 : 1;
	35352 : 1;
	35353 : 1;
	35354 : 1;
	35355 : 1;
	35356 : 1;
	35357 : 1;
	35358 : 1;
	35359 : 1;
	35360 : 1;
	35361 : 1;
	35362 : 1;
	35363 : 1;
	35364 : 1;
	35365 : 1;
	35366 : 1;
	35367 : 1;
	35368 : 1;
	35369 : 1;
	35370 : 1;
	35371 : 1;
	35372 : 1;
	35373 : 1;
	35374 : 1;
	35375 : 1;
	35376 : 1;
	35377 : 1;
	35378 : 1;
	35379 : 1;
	35380 : 1;
	35381 : 1;
	35382 : 1;
	35383 : 1;
	35384 : 1;
	35385 : 1;
	35386 : 1;
	35387 : 1;
	35388 : 1;
	35389 : 1;
	35390 : 1;
	35391 : 1;
	35392 : 1;
	35393 : 1;
	35394 : 1;
	35395 : 1;
	35396 : 1;
	35397 : 1;
	35398 : 1;
	35399 : 1;
	35400 : 1;
	35401 : 1;
	35402 : 1;
	35403 : 1;
	35404 : 1;
	35405 : 1;
	35406 : 1;
	35407 : 1;
	35408 : 1;
	35409 : 1;
	35410 : 1;
	35411 : 1;
	35412 : 1;
	35413 : 1;
	35414 : 1;
	35415 : 1;
	35416 : 1;
	35417 : 1;
	35418 : 1;
	35419 : 1;
	35420 : 1;
	35421 : 1;
	35422 : 1;
	35423 : 1;
	35424 : 1;
	35425 : 1;
	35426 : 1;
	35427 : 1;
	35428 : 1;
	35429 : 1;
	35430 : 1;
	35431 : 1;
	35432 : 1;
	35433 : 1;
	35434 : 1;
	35435 : 1;
	35436 : 1;
	35437 : 1;
	35438 : 1;
	35439 : 1;
	35440 : 1;
	35441 : 1;
	35442 : 1;
	35443 : 1;
	35444 : 1;
	35445 : 1;
	35446 : 1;
	35447 : 1;
	35448 : 1;
	35449 : 1;
	35450 : 1;
	35451 : 1;
	35452 : 1;
	35453 : 1;
	35454 : 1;
	35455 : 1;
	35456 : 1;
	35457 : 1;
	35458 : 1;
	35459 : 1;
	35460 : 1;
	35461 : 1;
	35462 : 1;
	35463 : 1;
	35464 : 1;
	35465 : 1;
	35466 : 1;
	35467 : 1;
	35468 : 1;
	35469 : 1;
	35470 : 1;
	35471 : 1;
	35472 : 1;
	35473 : 1;
	35474 : 1;
	35475 : 1;
	35476 : 1;
	35477 : 1;
	35478 : 1;
	35479 : 1;
	35480 : 1;
	35481 : 1;
	35482 : 1;
	35483 : 1;
	35484 : 1;
	35485 : 1;
	35486 : 1;
	35487 : 1;
	35488 : 1;
	35489 : 1;
	35490 : 1;
	35491 : 1;
	35492 : 1;
	35493 : 1;
	35494 : 1;
	35495 : 1;
	35496 : 1;
	35497 : 1;
	35498 : 1;
	35499 : 1;
	35500 : 1;
	35501 : 1;
	35502 : 1;
	35503 : 1;
	35504 : 1;
	35505 : 1;
	35506 : 1;
	35507 : 1;
	35508 : 1;
	35509 : 1;
	35510 : 1;
	35511 : 1;
	35512 : 1;
	35513 : 1;
	35514 : 1;
	35515 : 1;
	35516 : 1;
	35517 : 1;
	35518 : 1;
	35519 : 1;
	35520 : 1;
	35521 : 1;
	35522 : 1;
	35523 : 1;
	35524 : 1;
	35525 : 1;
	35526 : 1;
	35527 : 1;
	35528 : 1;
	35529 : 1;
	35530 : 1;
	35531 : 1;
	35532 : 1;
	35533 : 1;
	35534 : 1;
	35535 : 1;
	35536 : 1;
	35537 : 1;
	35538 : 1;
	35539 : 1;
	35540 : 1;
	35541 : 0;
	35542 : 0;
	35543 : 1;
	35544 : 1;
	35545 : 0;
	35546 : 1;
	35547 : 1;
	35548 : 1;
	35549 : 1;
	35550 : 1;
	35551 : 1;
	35552 : 1;
	35553 : 1;
	35554 : 1;
	35555 : 1;
	35556 : 0;
	35557 : 1;
	35558 : 1;
	35559 : 1;
	35560 : 1;
	35561 : 1;
	35562 : 1;
	35563 : 1;
	35564 : 1;
	35565 : 1;
	35566 : 1;
	35567 : 1;
	35568 : 1;
	35569 : 1;
	35570 : 1;
	35571 : 1;
	35572 : 0;
	35573 : 0;
	35574 : 1;
	35575 : 1;
	35576 : 0;
	35577 : 0;
	35578 : 0;
	35579 : 0;
	35580 : 1;
	35581 : 1;
	35582 : 1;
	35583 : 0;
	35584 : 1;
	35585 : 1;
	35586 : 1;
	35587 : 1;
	35588 : 1;
	35589 : 1;
	35590 : 0;
	35591 : 1;
	35592 : 1;
	35593 : 1;
	35594 : 1;
	35595 : 1;
	35596 : 1;
	35597 : 1;
	35598 : 1;
	35599 : 1;
	35600 : 1;
	35601 : 1;
	35602 : 1;
	35603 : 1;
	35604 : 1;
	35605 : 1;
	35606 : 1;
	35607 : 1;
	35608 : 1;
	35609 : 1;
	35610 : 1;
	35611 : 1;
	35612 : 1;
	35613 : 1;
	35614 : 1;
	35615 : 1;
	35616 : 1;
	35617 : 1;
	35618 : 1;
	35619 : 1;
	35620 : 1;
	35621 : 1;
	35622 : 1;
	35623 : 1;
	35624 : 1;
	35625 : 1;
	35626 : 1;
	35627 : 1;
	35628 : 1;
	35629 : 1;
	35630 : 1;
	35631 : 1;
	35632 : 1;
	35633 : 1;
	35634 : 1;
	35635 : 1;
	35636 : 1;
	35637 : 1;
	35638 : 1;
	35639 : 1;
	35640 : 1;
	35641 : 1;
	35642 : 1;
	35643 : 1;
	35644 : 1;
	35645 : 1;
	35646 : 1;
	35647 : 1;
	35648 : 1;
	35649 : 1;
	35650 : 1;
	35651 : 1;
	35652 : 1;
	35653 : 1;
	35654 : 1;
	35655 : 1;
	35656 : 1;
	35657 : 1;
	35658 : 1;
	35659 : 1;
	35660 : 1;
	35661 : 1;
	35662 : 1;
	35663 : 1;
	35664 : 1;
	35665 : 1;
	35666 : 1;
	35667 : 1;
	35668 : 1;
	35669 : 1;
	35670 : 1;
	35671 : 1;
	35672 : 1;
	35673 : 1;
	35674 : 1;
	35675 : 1;
	35676 : 1;
	35677 : 1;
	35678 : 1;
	35679 : 1;
	35680 : 1;
	35681 : 1;
	35682 : 1;
	35683 : 1;
	35684 : 1;
	35685 : 1;
	35686 : 1;
	35687 : 1;
	35688 : 1;
	35689 : 1;
	35690 : 1;
	35691 : 1;
	35692 : 1;
	35693 : 1;
	35694 : 1;
	35695 : 1;
	35696 : 1;
	35697 : 1;
	35698 : 1;
	35699 : 1;
	35700 : 1;
	35701 : 1;
	35702 : 1;
	35703 : 1;
	35704 : 1;
	35705 : 1;
	35706 : 1;
	35707 : 1;
	35708 : 1;
	35709 : 1;
	35710 : 1;
	35711 : 1;
	35712 : 1;
	35713 : 1;
	35714 : 1;
	35715 : 1;
	35716 : 1;
	35717 : 1;
	35718 : 1;
	35719 : 1;
	35720 : 1;
	35721 : 1;
	35722 : 1;
	35723 : 1;
	35724 : 1;
	35725 : 1;
	35726 : 1;
	35727 : 1;
	35728 : 1;
	35729 : 1;
	35730 : 1;
	35731 : 1;
	35732 : 1;
	35733 : 1;
	35734 : 1;
	35735 : 1;
	35736 : 1;
	35737 : 1;
	35738 : 1;
	35739 : 1;
	35740 : 1;
	35741 : 1;
	35742 : 1;
	35743 : 1;
	35744 : 1;
	35745 : 1;
	35746 : 1;
	35747 : 1;
	35748 : 1;
	35749 : 1;
	35750 : 1;
	35751 : 1;
	35752 : 1;
	35753 : 1;
	35754 : 1;
	35755 : 1;
	35756 : 1;
	35757 : 1;
	35758 : 1;
	35759 : 1;
	35760 : 1;
	35761 : 1;
	35762 : 1;
	35763 : 1;
	35764 : 1;
	35765 : 1;
	35766 : 1;
	35767 : 1;
	35768 : 1;
	35769 : 1;
	35770 : 1;
	35771 : 1;
	35772 : 1;
	35773 : 1;
	35774 : 1;
	35775 : 1;
	35776 : 1;
	35777 : 1;
	35778 : 1;
	35779 : 1;
	35780 : 1;
	35781 : 0;
	35782 : 0;
	35783 : 1;
	35784 : 1;
	35785 : 0;
	35786 : 1;
	35787 : 1;
	35788 : 1;
	35789 : 1;
	35790 : 1;
	35791 : 1;
	35792 : 1;
	35793 : 1;
	35794 : 1;
	35795 : 1;
	35796 : 0;
	35797 : 1;
	35798 : 1;
	35799 : 1;
	35800 : 1;
	35801 : 1;
	35802 : 1;
	35803 : 1;
	35804 : 1;
	35805 : 1;
	35806 : 1;
	35807 : 1;
	35808 : 1;
	35809 : 1;
	35810 : 1;
	35811 : 1;
	35812 : 0;
	35813 : 0;
	35814 : 1;
	35815 : 1;
	35816 : 0;
	35817 : 0;
	35818 : 1;
	35819 : 0;
	35820 : 1;
	35821 : 1;
	35822 : 1;
	35823 : 0;
	35824 : 0;
	35825 : 1;
	35826 : 1;
	35827 : 1;
	35828 : 1;
	35829 : 1;
	35830 : 0;
	35831 : 0;
	35832 : 1;
	35833 : 1;
	35834 : 1;
	35835 : 1;
	35836 : 1;
	35837 : 1;
	35838 : 1;
	35839 : 1;
	35840 : 1;
	35841 : 1;
	35842 : 1;
	35843 : 1;
	35844 : 1;
	35845 : 1;
	35846 : 1;
	35847 : 1;
	35848 : 1;
	35849 : 1;
	35850 : 1;
	35851 : 1;
	35852 : 1;
	35853 : 1;
	35854 : 1;
	35855 : 1;
	35856 : 1;
	35857 : 1;
	35858 : 1;
	35859 : 1;
	35860 : 1;
	35861 : 1;
	35862 : 1;
	35863 : 1;
	35864 : 1;
	35865 : 1;
	35866 : 1;
	35867 : 1;
	35868 : 1;
	35869 : 1;
	35870 : 1;
	35871 : 1;
	35872 : 1;
	35873 : 1;
	35874 : 1;
	35875 : 1;
	35876 : 1;
	35877 : 1;
	35878 : 1;
	35879 : 1;
	35880 : 1;
	35881 : 1;
	35882 : 1;
	35883 : 1;
	35884 : 1;
	35885 : 1;
	35886 : 1;
	35887 : 1;
	35888 : 1;
	35889 : 1;
	35890 : 1;
	35891 : 1;
	35892 : 1;
	35893 : 1;
	35894 : 1;
	35895 : 1;
	35896 : 1;
	35897 : 1;
	35898 : 1;
	35899 : 1;
	35900 : 1;
	35901 : 1;
	35902 : 1;
	35903 : 1;
	35904 : 1;
	35905 : 1;
	35906 : 1;
	35907 : 1;
	35908 : 1;
	35909 : 1;
	35910 : 1;
	35911 : 1;
	35912 : 1;
	35913 : 1;
	35914 : 1;
	35915 : 1;
	35916 : 1;
	35917 : 1;
	35918 : 1;
	35919 : 1;
	35920 : 1;
	35921 : 1;
	35922 : 1;
	35923 : 1;
	35924 : 1;
	35925 : 1;
	35926 : 0;
	35927 : 0;
	35928 : 0;
	35929 : 0;
	35930 : 1;
	35931 : 1;
	35932 : 1;
	35933 : 1;
	35934 : 1;
	35935 : 0;
	35936 : 1;
	35937 : 1;
	35938 : 1;
	35939 : 1;
	35940 : 1;
	35941 : 1;
	35942 : 1;
	35943 : 1;
	35944 : 1;
	35945 : 1;
	35946 : 1;
	35947 : 1;
	35948 : 1;
	35949 : 0;
	35950 : 1;
	35951 : 1;
	35952 : 1;
	35953 : 1;
	35954 : 1;
	35955 : 1;
	35956 : 1;
	35957 : 1;
	35958 : 1;
	35959 : 1;
	35960 : 1;
	35961 : 1;
	35962 : 1;
	35963 : 0;
	35964 : 0;
	35965 : 1;
	35966 : 1;
	35967 : 1;
	35968 : 1;
	35969 : 1;
	35970 : 1;
	35971 : 1;
	35972 : 1;
	35973 : 1;
	35974 : 1;
	35975 : 1;
	35976 : 1;
	35977 : 1;
	35978 : 1;
	35979 : 1;
	35980 : 1;
	35981 : 1;
	35982 : 1;
	35983 : 1;
	35984 : 1;
	35985 : 1;
	35986 : 1;
	35987 : 1;
	35988 : 1;
	35989 : 1;
	35990 : 1;
	35991 : 1;
	35992 : 1;
	35993 : 1;
	35994 : 1;
	35995 : 1;
	35996 : 1;
	35997 : 1;
	35998 : 1;
	35999 : 1;
	36000 : 1;
	36001 : 1;
	36002 : 1;
	36003 : 1;
	36004 : 1;
	36005 : 0;
	36006 : 0;
	36007 : 0;
	36008 : 1;
	36009 : 0;
	36010 : 0;
	36011 : 0;
	36012 : 0;
	36013 : 1;
	36014 : 0;
	36015 : 0;
	36016 : 0;
	36017 : 1;
	36018 : 1;
	36019 : 0;
	36020 : 0;
	36021 : 0;
	36022 : 0;
	36023 : 1;
	36024 : 1;
	36025 : 0;
	36026 : 1;
	36027 : 0;
	36028 : 1;
	36029 : 0;
	36030 : 1;
	36031 : 1;
	36032 : 0;
	36033 : 0;
	36034 : 0;
	36035 : 1;
	36036 : 0;
	36037 : 1;
	36038 : 0;
	36039 : 0;
	36040 : 1;
	36041 : 1;
	36042 : 0;
	36043 : 0;
	36044 : 0;
	36045 : 0;
	36046 : 1;
	36047 : 1;
	36048 : 1;
	36049 : 1;
	36050 : 0;
	36051 : 0;
	36052 : 0;
	36053 : 1;
	36054 : 0;
	36055 : 0;
	36056 : 0;
	36057 : 0;
	36058 : 1;
	36059 : 0;
	36060 : 1;
	36061 : 1;
	36062 : 1;
	36063 : 1;
	36064 : 1;
	36065 : 0;
	36066 : 0;
	36067 : 0;
	36068 : 0;
	36069 : 1;
	36070 : 1;
	36071 : 1;
	36072 : 1;
	36073 : 1;
	36074 : 1;
	36075 : 1;
	36076 : 1;
	36077 : 1;
	36078 : 1;
	36079 : 1;
	36080 : 1;
	36081 : 1;
	36082 : 1;
	36083 : 1;
	36084 : 1;
	36085 : 1;
	36086 : 1;
	36087 : 1;
	36088 : 1;
	36089 : 1;
	36090 : 1;
	36091 : 1;
	36092 : 1;
	36093 : 1;
	36094 : 1;
	36095 : 1;
	36096 : 1;
	36097 : 1;
	36098 : 1;
	36099 : 1;
	36100 : 1;
	36101 : 1;
	36102 : 1;
	36103 : 1;
	36104 : 1;
	36105 : 1;
	36106 : 1;
	36107 : 1;
	36108 : 1;
	36109 : 1;
	36110 : 1;
	36111 : 1;
	36112 : 1;
	36113 : 1;
	36114 : 1;
	36115 : 1;
	36116 : 1;
	36117 : 1;
	36118 : 1;
	36119 : 1;
	36120 : 1;
	36121 : 1;
	36122 : 1;
	36123 : 1;
	36124 : 1;
	36125 : 1;
	36126 : 1;
	36127 : 1;
	36128 : 1;
	36129 : 1;
	36130 : 1;
	36131 : 1;
	36132 : 1;
	36133 : 1;
	36134 : 1;
	36135 : 1;
	36136 : 1;
	36137 : 1;
	36138 : 1;
	36139 : 1;
	36140 : 1;
	36141 : 1;
	36142 : 1;
	36143 : 1;
	36144 : 1;
	36145 : 1;
	36146 : 1;
	36147 : 1;
	36148 : 1;
	36149 : 1;
	36150 : 1;
	36151 : 1;
	36152 : 1;
	36153 : 1;
	36154 : 1;
	36155 : 1;
	36156 : 1;
	36157 : 1;
	36158 : 1;
	36159 : 1;
	36160 : 1;
	36161 : 1;
	36162 : 1;
	36163 : 1;
	36164 : 1;
	36165 : 1;
	36166 : 0;
	36167 : 1;
	36168 : 1;
	36169 : 1;
	36170 : 1;
	36171 : 1;
	36172 : 1;
	36173 : 1;
	36174 : 1;
	36175 : 0;
	36176 : 1;
	36177 : 1;
	36178 : 1;
	36179 : 1;
	36180 : 1;
	36181 : 1;
	36182 : 1;
	36183 : 1;
	36184 : 1;
	36185 : 1;
	36186 : 1;
	36187 : 1;
	36188 : 1;
	36189 : 0;
	36190 : 1;
	36191 : 1;
	36192 : 1;
	36193 : 1;
	36194 : 1;
	36195 : 1;
	36196 : 1;
	36197 : 1;
	36198 : 1;
	36199 : 1;
	36200 : 1;
	36201 : 1;
	36202 : 1;
	36203 : 1;
	36204 : 0;
	36205 : 1;
	36206 : 1;
	36207 : 1;
	36208 : 1;
	36209 : 1;
	36210 : 1;
	36211 : 1;
	36212 : 1;
	36213 : 1;
	36214 : 1;
	36215 : 1;
	36216 : 1;
	36217 : 1;
	36218 : 1;
	36219 : 1;
	36220 : 1;
	36221 : 1;
	36222 : 1;
	36223 : 1;
	36224 : 1;
	36225 : 1;
	36226 : 1;
	36227 : 1;
	36228 : 1;
	36229 : 1;
	36230 : 1;
	36231 : 1;
	36232 : 1;
	36233 : 1;
	36234 : 1;
	36235 : 1;
	36236 : 1;
	36237 : 1;
	36238 : 1;
	36239 : 1;
	36240 : 1;
	36241 : 1;
	36242 : 1;
	36243 : 1;
	36244 : 0;
	36245 : 1;
	36246 : 1;
	36247 : 0;
	36248 : 1;
	36249 : 0;
	36250 : 1;
	36251 : 1;
	36252 : 0;
	36253 : 1;
	36254 : 0;
	36255 : 1;
	36256 : 1;
	36257 : 0;
	36258 : 0;
	36259 : 1;
	36260 : 1;
	36261 : 0;
	36262 : 0;
	36263 : 1;
	36264 : 1;
	36265 : 0;
	36266 : 1;
	36267 : 0;
	36268 : 1;
	36269 : 0;
	36270 : 1;
	36271 : 1;
	36272 : 0;
	36273 : 1;
	36274 : 1;
	36275 : 0;
	36276 : 0;
	36277 : 0;
	36278 : 0;
	36279 : 1;
	36280 : 1;
	36281 : 1;
	36282 : 0;
	36283 : 0;
	36284 : 1;
	36285 : 1;
	36286 : 0;
	36287 : 1;
	36288 : 1;
	36289 : 1;
	36290 : 1;
	36291 : 1;
	36292 : 0;
	36293 : 1;
	36294 : 1;
	36295 : 1;
	36296 : 0;
	36297 : 0;
	36298 : 1;
	36299 : 0;
	36300 : 1;
	36301 : 1;
	36302 : 1;
	36303 : 1;
	36304 : 1;
	36305 : 1;
	36306 : 1;
	36307 : 1;
	36308 : 1;
	36309 : 1;
	36310 : 1;
	36311 : 1;
	36312 : 1;
	36313 : 1;
	36314 : 1;
	36315 : 1;
	36316 : 1;
	36317 : 1;
	36318 : 1;
	36319 : 1;
	36320 : 1;
	36321 : 1;
	36322 : 1;
	36323 : 1;
	36324 : 1;
	36325 : 1;
	36326 : 1;
	36327 : 1;
	36328 : 1;
	36329 : 1;
	36330 : 1;
	36331 : 1;
	36332 : 1;
	36333 : 1;
	36334 : 1;
	36335 : 1;
	36336 : 1;
	36337 : 1;
	36338 : 1;
	36339 : 1;
	36340 : 1;
	36341 : 1;
	36342 : 1;
	36343 : 1;
	36344 : 1;
	36345 : 1;
	36346 : 1;
	36347 : 1;
	36348 : 1;
	36349 : 1;
	36350 : 1;
	36351 : 1;
	36352 : 1;
	36353 : 1;
	36354 : 1;
	36355 : 1;
	36356 : 1;
	36357 : 1;
	36358 : 1;
	36359 : 1;
	36360 : 1;
	36361 : 1;
	36362 : 1;
	36363 : 1;
	36364 : 1;
	36365 : 1;
	36366 : 1;
	36367 : 1;
	36368 : 1;
	36369 : 1;
	36370 : 1;
	36371 : 1;
	36372 : 1;
	36373 : 1;
	36374 : 1;
	36375 : 1;
	36376 : 1;
	36377 : 1;
	36378 : 1;
	36379 : 1;
	36380 : 1;
	36381 : 1;
	36382 : 1;
	36383 : 0;
	36384 : 0;
	36385 : 0;
	36386 : 0;
	36387 : 1;
	36388 : 0;
	36389 : 0;
	36390 : 0;
	36391 : 1;
	36392 : 0;
	36393 : 0;
	36394 : 0;
	36395 : 1;
	36396 : 0;
	36397 : 0;
	36398 : 0;
	36399 : 0;
	36400 : 0;
	36401 : 0;
	36402 : 0;
	36403 : 0;
	36404 : 1;
	36405 : 1;
	36406 : 0;
	36407 : 0;
	36408 : 0;
	36409 : 1;
	36410 : 0;
	36411 : 0;
	36412 : 0;
	36413 : 1;
	36414 : 0;
	36415 : 0;
	36416 : 0;
	36417 : 0;
	36418 : 1;
	36419 : 0;
	36420 : 0;
	36421 : 0;
	36422 : 1;
	36423 : 0;
	36424 : 0;
	36425 : 0;
	36426 : 1;
	36427 : 1;
	36428 : 0;
	36429 : 0;
	36430 : 0;
	36431 : 0;
	36432 : 1;
	36433 : 0;
	36434 : 0;
	36435 : 0;
	36436 : 1;
	36437 : 1;
	36438 : 0;
	36439 : 0;
	36440 : 0;
	36441 : 0;
	36442 : 1;
	36443 : 1;
	36444 : 0;
	36445 : 1;
	36446 : 0;
	36447 : 0;
	36448 : 0;
	36449 : 0;
	36450 : 0;
	36451 : 1;
	36452 : 1;
	36453 : 0;
	36454 : 1;
	36455 : 1;
	36456 : 1;
	36457 : 0;
	36458 : 0;
	36459 : 0;
	36460 : 0;
	36461 : 1;
	36462 : 0;
	36463 : 0;
	36464 : 0;
	36465 : 1;
	36466 : 0;
	36467 : 0;
	36468 : 0;
	36469 : 0;
	36470 : 0;
	36471 : 1;
	36472 : 0;
	36473 : 0;
	36474 : 0;
	36475 : 1;
	36476 : 1;
	36477 : 1;
	36478 : 1;
	36479 : 1;
	36480 : 1;
	36481 : 1;
	36482 : 1;
	36483 : 1;
	36484 : 0;
	36485 : 1;
	36486 : 1;
	36487 : 0;
	36488 : 1;
	36489 : 0;
	36490 : 1;
	36491 : 1;
	36492 : 0;
	36493 : 1;
	36494 : 0;
	36495 : 1;
	36496 : 1;
	36497 : 0;
	36498 : 0;
	36499 : 1;
	36500 : 1;
	36501 : 0;
	36502 : 0;
	36503 : 1;
	36504 : 1;
	36505 : 0;
	36506 : 1;
	36507 : 0;
	36508 : 1;
	36509 : 0;
	36510 : 1;
	36511 : 1;
	36512 : 0;
	36513 : 1;
	36514 : 1;
	36515 : 0;
	36516 : 0;
	36517 : 0;
	36518 : 1;
	36519 : 1;
	36520 : 1;
	36521 : 1;
	36522 : 0;
	36523 : 0;
	36524 : 1;
	36525 : 1;
	36526 : 0;
	36527 : 1;
	36528 : 1;
	36529 : 1;
	36530 : 1;
	36531 : 1;
	36532 : 0;
	36533 : 1;
	36534 : 1;
	36535 : 1;
	36536 : 0;
	36537 : 0;
	36538 : 1;
	36539 : 0;
	36540 : 1;
	36541 : 1;
	36542 : 1;
	36543 : 0;
	36544 : 0;
	36545 : 1;
	36546 : 1;
	36547 : 1;
	36548 : 1;
	36549 : 1;
	36550 : 0;
	36551 : 0;
	36552 : 1;
	36553 : 1;
	36554 : 1;
	36555 : 1;
	36556 : 1;
	36557 : 1;
	36558 : 1;
	36559 : 1;
	36560 : 1;
	36561 : 1;
	36562 : 1;
	36563 : 1;
	36564 : 1;
	36565 : 1;
	36566 : 1;
	36567 : 1;
	36568 : 1;
	36569 : 1;
	36570 : 1;
	36571 : 1;
	36572 : 1;
	36573 : 1;
	36574 : 1;
	36575 : 1;
	36576 : 1;
	36577 : 1;
	36578 : 1;
	36579 : 1;
	36580 : 1;
	36581 : 1;
	36582 : 1;
	36583 : 1;
	36584 : 1;
	36585 : 1;
	36586 : 1;
	36587 : 1;
	36588 : 1;
	36589 : 1;
	36590 : 1;
	36591 : 1;
	36592 : 1;
	36593 : 1;
	36594 : 1;
	36595 : 1;
	36596 : 1;
	36597 : 1;
	36598 : 1;
	36599 : 1;
	36600 : 1;
	36601 : 1;
	36602 : 1;
	36603 : 1;
	36604 : 1;
	36605 : 1;
	36606 : 1;
	36607 : 1;
	36608 : 1;
	36609 : 1;
	36610 : 1;
	36611 : 1;
	36612 : 1;
	36613 : 1;
	36614 : 1;
	36615 : 1;
	36616 : 1;
	36617 : 1;
	36618 : 1;
	36619 : 1;
	36620 : 1;
	36621 : 1;
	36622 : 1;
	36623 : 0;
	36624 : 1;
	36625 : 1;
	36626 : 0;
	36627 : 1;
	36628 : 0;
	36629 : 1;
	36630 : 1;
	36631 : 1;
	36632 : 0;
	36633 : 0;
	36634 : 0;
	36635 : 0;
	36636 : 0;
	36637 : 0;
	36638 : 0;
	36639 : 1;
	36640 : 0;
	36641 : 0;
	36642 : 1;
	36643 : 1;
	36644 : 1;
	36645 : 1;
	36646 : 0;
	36647 : 1;
	36648 : 1;
	36649 : 1;
	36650 : 0;
	36651 : 1;
	36652 : 1;
	36653 : 0;
	36654 : 1;
	36655 : 0;
	36656 : 1;
	36657 : 1;
	36658 : 0;
	36659 : 0;
	36660 : 0;
	36661 : 0;
	36662 : 1;
	36663 : 0;
	36664 : 0;
	36665 : 1;
	36666 : 1;
	36667 : 1;
	36668 : 1;
	36669 : 0;
	36670 : 1;
	36671 : 1;
	36672 : 0;
	36673 : 1;
	36674 : 1;
	36675 : 0;
	36676 : 1;
	36677 : 1;
	36678 : 0;
	36679 : 1;
	36680 : 1;
	36681 : 0;
	36682 : 0;
	36683 : 1;
	36684 : 0;
	36685 : 0;
	36686 : 1;
	36687 : 1;
	36688 : 0;
	36689 : 0;
	36690 : 0;
	36691 : 1;
	36692 : 1;
	36693 : 0;
	36694 : 1;
	36695 : 1;
	36696 : 0;
	36697 : 1;
	36698 : 1;
	36699 : 0;
	36700 : 0;
	36701 : 0;
	36702 : 1;
	36703 : 1;
	36704 : 0;
	36705 : 1;
	36706 : 0;
	36707 : 1;
	36708 : 1;
	36709 : 0;
	36710 : 0;
	36711 : 1;
	36712 : 0;
	36713 : 1;
	36714 : 0;
	36715 : 0;
	36716 : 1;
	36717 : 1;
	36718 : 1;
	36719 : 1;
	36720 : 1;
	36721 : 1;
	36722 : 1;
	36723 : 1;
	36724 : 1;
	36725 : 0;
	36726 : 0;
	36727 : 0;
	36728 : 1;
	36729 : 0;
	36730 : 0;
	36731 : 0;
	36732 : 0;
	36733 : 1;
	36734 : 0;
	36735 : 0;
	36736 : 0;
	36737 : 1;
	36738 : 1;
	36739 : 0;
	36740 : 0;
	36741 : 0;
	36742 : 0;
	36743 : 1;
	36744 : 1;
	36745 : 0;
	36746 : 1;
	36747 : 0;
	36748 : 0;
	36749 : 0;
	36750 : 0;
	36751 : 1;
	36752 : 0;
	36753 : 0;
	36754 : 0;
	36755 : 1;
	36756 : 0;
	36757 : 1;
	36758 : 0;
	36759 : 0;
	36760 : 1;
	36761 : 1;
	36762 : 0;
	36763 : 0;
	36764 : 1;
	36765 : 1;
	36766 : 0;
	36767 : 1;
	36768 : 1;
	36769 : 0;
	36770 : 0;
	36771 : 0;
	36772 : 1;
	36773 : 1;
	36774 : 0;
	36775 : 0;
	36776 : 0;
	36777 : 1;
	36778 : 0;
	36779 : 0;
	36780 : 0;
	36781 : 1;
	36782 : 1;
	36783 : 0;
	36784 : 0;
	36785 : 1;
	36786 : 1;
	36787 : 1;
	36788 : 1;
	36789 : 1;
	36790 : 0;
	36791 : 0;
	36792 : 1;
	36793 : 1;
	36794 : 1;
	36795 : 1;
	36796 : 1;
	36797 : 1;
	36798 : 1;
	36799 : 1;
	36800 : 1;
	36801 : 1;
	36802 : 1;
	36803 : 1;
	36804 : 1;
	36805 : 1;
	36806 : 1;
	36807 : 1;
	36808 : 1;
	36809 : 1;
	36810 : 1;
	36811 : 1;
	36812 : 1;
	36813 : 1;
	36814 : 1;
	36815 : 1;
	36816 : 1;
	36817 : 1;
	36818 : 1;
	36819 : 1;
	36820 : 1;
	36821 : 1;
	36822 : 1;
	36823 : 1;
	36824 : 1;
	36825 : 1;
	36826 : 1;
	36827 : 1;
	36828 : 1;
	36829 : 1;
	36830 : 1;
	36831 : 1;
	36832 : 1;
	36833 : 1;
	36834 : 1;
	36835 : 1;
	36836 : 1;
	36837 : 1;
	36838 : 1;
	36839 : 1;
	36840 : 1;
	36841 : 1;
	36842 : 1;
	36843 : 1;
	36844 : 1;
	36845 : 1;
	36846 : 1;
	36847 : 1;
	36848 : 1;
	36849 : 1;
	36850 : 1;
	36851 : 1;
	36852 : 1;
	36853 : 1;
	36854 : 1;
	36855 : 1;
	36856 : 1;
	36857 : 1;
	36858 : 1;
	36859 : 1;
	36860 : 1;
	36861 : 1;
	36862 : 1;
	36863 : 0;
	36864 : 1;
	36865 : 1;
	36866 : 0;
	36867 : 1;
	36868 : 0;
	36869 : 1;
	36870 : 1;
	36871 : 1;
	36872 : 0;
	36873 : 0;
	36874 : 0;
	36875 : 0;
	36876 : 1;
	36877 : 0;
	36878 : 0;
	36879 : 0;
	36880 : 1;
	36881 : 0;
	36882 : 0;
	36883 : 1;
	36884 : 1;
	36885 : 1;
	36886 : 0;
	36887 : 1;
	36888 : 1;
	36889 : 1;
	36890 : 0;
	36891 : 1;
	36892 : 1;
	36893 : 0;
	36894 : 1;
	36895 : 0;
	36896 : 1;
	36897 : 1;
	36898 : 0;
	36899 : 0;
	36900 : 0;
	36901 : 0;
	36902 : 1;
	36903 : 0;
	36904 : 1;
	36905 : 1;
	36906 : 1;
	36907 : 1;
	36908 : 1;
	36909 : 0;
	36910 : 1;
	36911 : 1;
	36912 : 0;
	36913 : 1;
	36914 : 1;
	36915 : 0;
	36916 : 1;
	36917 : 1;
	36918 : 0;
	36919 : 1;
	36920 : 1;
	36921 : 0;
	36922 : 0;
	36923 : 1;
	36924 : 0;
	36925 : 0;
	36926 : 1;
	36927 : 1;
	36928 : 0;
	36929 : 0;
	36930 : 0;
	36931 : 1;
	36932 : 1;
	36933 : 0;
	36934 : 1;
	36935 : 1;
	36936 : 0;
	36937 : 1;
	36938 : 1;
	36939 : 0;
	36940 : 0;
	36941 : 0;
	36942 : 1;
	36943 : 1;
	36944 : 0;
	36945 : 1;
	36946 : 0;
	36947 : 1;
	36948 : 0;
	36949 : 0;
	36950 : 0;
	36951 : 1;
	36952 : 0;
	36953 : 1;
	36954 : 0;
	36955 : 0;
	36956 : 1;
	36957 : 1;
	36958 : 1;
	36959 : 1;
	36960 : 1;
	36961 : 1;
	36962 : 1;
	36963 : 1;
	36964 : 1;
	36965 : 0;
	36966 : 0;
	36967 : 0;
	36968 : 1;
	36969 : 1;
	36970 : 1;
	36971 : 1;
	36972 : 1;
	36973 : 1;
	36974 : 1;
	36975 : 1;
	36976 : 1;
	36977 : 1;
	36978 : 1;
	36979 : 1;
	36980 : 1;
	36981 : 1;
	36982 : 1;
	36983 : 1;
	36984 : 1;
	36985 : 1;
	36986 : 1;
	36987 : 1;
	36988 : 1;
	36989 : 1;
	36990 : 1;
	36991 : 1;
	36992 : 1;
	36993 : 1;
	36994 : 1;
	36995 : 1;
	36996 : 1;
	36997 : 1;
	36998 : 1;
	36999 : 1;
	37000 : 1;
	37001 : 1;
	37002 : 1;
	37003 : 1;
	37004 : 1;
	37005 : 1;
	37006 : 1;
	37007 : 1;
	37008 : 1;
	37009 : 1;
	37010 : 1;
	37011 : 1;
	37012 : 1;
	37013 : 1;
	37014 : 1;
	37015 : 1;
	37016 : 1;
	37017 : 1;
	37018 : 1;
	37019 : 1;
	37020 : 1;
	37021 : 1;
	37022 : 1;
	37023 : 0;
	37024 : 1;
	37025 : 1;
	37026 : 1;
	37027 : 1;
	37028 : 1;
	37029 : 1;
	37030 : 0;
	37031 : 1;
	37032 : 1;
	37033 : 1;
	37034 : 1;
	37035 : 1;
	37036 : 1;
	37037 : 1;
	37038 : 1;
	37039 : 1;
	37040 : 1;
	37041 : 1;
	37042 : 1;
	37043 : 1;
	37044 : 1;
	37045 : 1;
	37046 : 1;
	37047 : 1;
	37048 : 1;
	37049 : 1;
	37050 : 1;
	37051 : 1;
	37052 : 1;
	37053 : 1;
	37054 : 1;
	37055 : 1;
	37056 : 1;
	37057 : 1;
	37058 : 1;
	37059 : 1;
	37060 : 1;
	37061 : 1;
	37062 : 1;
	37063 : 1;
	37064 : 1;
	37065 : 1;
	37066 : 1;
	37067 : 1;
	37068 : 1;
	37069 : 1;
	37070 : 1;
	37071 : 1;
	37072 : 1;
	37073 : 1;
	37074 : 1;
	37075 : 1;
	37076 : 1;
	37077 : 1;
	37078 : 1;
	37079 : 1;
	37080 : 1;
	37081 : 1;
	37082 : 1;
	37083 : 1;
	37084 : 1;
	37085 : 1;
	37086 : 1;
	37087 : 1;
	37088 : 1;
	37089 : 1;
	37090 : 1;
	37091 : 1;
	37092 : 1;
	37093 : 1;
	37094 : 1;
	37095 : 1;
	37096 : 1;
	37097 : 1;
	37098 : 1;
	37099 : 1;
	37100 : 1;
	37101 : 1;
	37102 : 1;
	37103 : 0;
	37104 : 0;
	37105 : 0;
	37106 : 0;
	37107 : 1;
	37108 : 0;
	37109 : 1;
	37110 : 1;
	37111 : 1;
	37112 : 0;
	37113 : 0;
	37114 : 0;
	37115 : 0;
	37116 : 0;
	37117 : 0;
	37118 : 0;
	37119 : 0;
	37120 : 0;
	37121 : 0;
	37122 : 0;
	37123 : 0;
	37124 : 1;
	37125 : 1;
	37126 : 0;
	37127 : 0;
	37128 : 0;
	37129 : 0;
	37130 : 0;
	37131 : 1;
	37132 : 1;
	37133 : 0;
	37134 : 1;
	37135 : 0;
	37136 : 0;
	37137 : 0;
	37138 : 1;
	37139 : 0;
	37140 : 0;
	37141 : 0;
	37142 : 1;
	37143 : 0;
	37144 : 1;
	37145 : 1;
	37146 : 1;
	37147 : 1;
	37148 : 1;
	37149 : 0;
	37150 : 0;
	37151 : 0;
	37152 : 1;
	37153 : 0;
	37154 : 0;
	37155 : 0;
	37156 : 1;
	37157 : 1;
	37158 : 0;
	37159 : 0;
	37160 : 0;
	37161 : 0;
	37162 : 1;
	37163 : 1;
	37164 : 0;
	37165 : 1;
	37166 : 0;
	37167 : 0;
	37168 : 0;
	37169 : 0;
	37170 : 1;
	37171 : 0;
	37172 : 0;
	37173 : 0;
	37174 : 1;
	37175 : 1;
	37176 : 1;
	37177 : 0;
	37178 : 0;
	37179 : 0;
	37180 : 0;
	37181 : 1;
	37182 : 0;
	37183 : 0;
	37184 : 0;
	37185 : 1;
	37186 : 0;
	37187 : 0;
	37188 : 0;
	37189 : 0;
	37190 : 0;
	37191 : 1;
	37192 : 0;
	37193 : 1;
	37194 : 0;
	37195 : 0;
	37196 : 1;
	37197 : 1;
	37198 : 1;
	37199 : 1;
	37200 : 1;
	37201 : 1;
	37202 : 1;
	37203 : 1;
	37204 : 1;
	37205 : 0;
	37206 : 0;
	37207 : 1;
	37208 : 1;
	37209 : 1;
	37210 : 1;
	37211 : 1;
	37212 : 1;
	37213 : 1;
	37214 : 1;
	37215 : 1;
	37216 : 1;
	37217 : 1;
	37218 : 1;
	37219 : 1;
	37220 : 1;
	37221 : 1;
	37222 : 1;
	37223 : 1;
	37224 : 1;
	37225 : 1;
	37226 : 1;
	37227 : 1;
	37228 : 1;
	37229 : 1;
	37230 : 1;
	37231 : 1;
	37232 : 1;
	37233 : 1;
	37234 : 1;
	37235 : 1;
	37236 : 1;
	37237 : 1;
	37238 : 1;
	37239 : 1;
	37240 : 1;
	37241 : 1;
	37242 : 1;
	37243 : 1;
	37244 : 1;
	37245 : 1;
	37246 : 1;
	37247 : 1;
	37248 : 1;
	37249 : 1;
	37250 : 1;
	37251 : 1;
	37252 : 1;
	37253 : 1;
	37254 : 1;
	37255 : 1;
	37256 : 1;
	37257 : 1;
	37258 : 1;
	37259 : 1;
	37260 : 1;
	37261 : 1;
	37262 : 1;
	37263 : 1;
	37264 : 1;
	37265 : 1;
	37266 : 1;
	37267 : 1;
	37268 : 1;
	37269 : 1;
	37270 : 1;
	37271 : 1;
	37272 : 1;
	37273 : 1;
	37274 : 1;
	37275 : 1;
	37276 : 1;
	37277 : 1;
	37278 : 1;
	37279 : 1;
	37280 : 1;
	37281 : 1;
	37282 : 1;
	37283 : 1;
	37284 : 1;
	37285 : 1;
	37286 : 1;
	37287 : 1;
	37288 : 1;
	37289 : 1;
	37290 : 1;
	37291 : 1;
	37292 : 1;
	37293 : 1;
	37294 : 1;
	37295 : 1;
	37296 : 1;
	37297 : 1;
	37298 : 1;
	37299 : 1;
	37300 : 1;
	37301 : 1;
	37302 : 1;
	37303 : 1;
	37304 : 1;
	37305 : 1;
	37306 : 1;
	37307 : 1;
	37308 : 1;
	37309 : 1;
	37310 : 1;
	37311 : 1;
	37312 : 1;
	37313 : 1;
	37314 : 1;
	37315 : 1;
	37316 : 1;
	37317 : 1;
	37318 : 1;
	37319 : 1;
	37320 : 1;
	37321 : 1;
	37322 : 1;
	37323 : 1;
	37324 : 1;
	37325 : 1;
	37326 : 1;
	37327 : 1;
	37328 : 1;
	37329 : 1;
	37330 : 1;
	37331 : 1;
	37332 : 1;
	37333 : 1;
	37334 : 1;
	37335 : 1;
	37336 : 1;
	37337 : 1;
	37338 : 1;
	37339 : 1;
	37340 : 1;
	37341 : 1;
	37342 : 1;
	37343 : 0;
	37344 : 1;
	37345 : 1;
	37346 : 1;
	37347 : 1;
	37348 : 1;
	37349 : 1;
	37350 : 1;
	37351 : 1;
	37352 : 1;
	37353 : 1;
	37354 : 1;
	37355 : 1;
	37356 : 1;
	37357 : 1;
	37358 : 1;
	37359 : 1;
	37360 : 1;
	37361 : 1;
	37362 : 1;
	37363 : 1;
	37364 : 1;
	37365 : 1;
	37366 : 1;
	37367 : 1;
	37368 : 1;
	37369 : 1;
	37370 : 1;
	37371 : 1;
	37372 : 1;
	37373 : 1;
	37374 : 1;
	37375 : 1;
	37376 : 1;
	37377 : 1;
	37378 : 1;
	37379 : 1;
	37380 : 1;
	37381 : 1;
	37382 : 1;
	37383 : 1;
	37384 : 1;
	37385 : 1;
	37386 : 1;
	37387 : 1;
	37388 : 1;
	37389 : 1;
	37390 : 1;
	37391 : 1;
	37392 : 1;
	37393 : 1;
	37394 : 1;
	37395 : 1;
	37396 : 1;
	37397 : 1;
	37398 : 0;
	37399 : 1;
	37400 : 1;
	37401 : 1;
	37402 : 1;
	37403 : 1;
	37404 : 1;
	37405 : 1;
	37406 : 1;
	37407 : 1;
	37408 : 1;
	37409 : 1;
	37410 : 1;
	37411 : 0;
	37412 : 0;
	37413 : 0;
	37414 : 1;
	37415 : 1;
	37416 : 1;
	37417 : 1;
	37418 : 1;
	37419 : 1;
	37420 : 1;
	37421 : 1;
	37422 : 0;
	37423 : 0;
	37424 : 0;
	37425 : 1;
	37426 : 1;
	37427 : 1;
	37428 : 1;
	37429 : 1;
	37430 : 1;
	37431 : 1;
	37432 : 1;
	37433 : 1;
	37434 : 1;
	37435 : 1;
	37436 : 1;
	37437 : 1;
	37438 : 1;
	37439 : 1;
	37440 : 1;
	37441 : 1;
	37442 : 1;
	37443 : 1;
	37444 : 1;
	37445 : 1;
	37446 : 1;
	37447 : 1;
	37448 : 1;
	37449 : 1;
	37450 : 1;
	37451 : 1;
	37452 : 1;
	37453 : 1;
	37454 : 1;
	37455 : 1;
	37456 : 1;
	37457 : 1;
	37458 : 1;
	37459 : 1;
	37460 : 1;
	37461 : 1;
	37462 : 1;
	37463 : 1;
	37464 : 1;
	37465 : 1;
	37466 : 1;
	37467 : 1;
	37468 : 1;
	37469 : 1;
	37470 : 1;
	37471 : 1;
	37472 : 1;
	37473 : 1;
	37474 : 1;
	37475 : 1;
	37476 : 1;
	37477 : 1;
	37478 : 1;
	37479 : 1;
	37480 : 1;
	37481 : 1;
	37482 : 1;
	37483 : 1;
	37484 : 1;
	37485 : 1;
	37486 : 1;
	37487 : 1;
	37488 : 1;
	37489 : 1;
	37490 : 1;
	37491 : 1;
	37492 : 1;
	37493 : 1;
	37494 : 1;
	37495 : 1;
	37496 : 1;
	37497 : 1;
	37498 : 1;
	37499 : 1;
	37500 : 1;
	37501 : 1;
	37502 : 1;
	37503 : 1;
	37504 : 1;
	37505 : 1;
	37506 : 1;
	37507 : 1;
	37508 : 1;
	37509 : 1;
	37510 : 1;
	37511 : 1;
	37512 : 1;
	37513 : 1;
	37514 : 1;
	37515 : 1;
	37516 : 1;
	37517 : 1;
	37518 : 1;
	37519 : 1;
	37520 : 1;
	37521 : 1;
	37522 : 1;
	37523 : 1;
	37524 : 1;
	37525 : 1;
	37526 : 1;
	37527 : 1;
	37528 : 1;
	37529 : 1;
	37530 : 1;
	37531 : 1;
	37532 : 1;
	37533 : 1;
	37534 : 1;
	37535 : 1;
	37536 : 1;
	37537 : 1;
	37538 : 1;
	37539 : 1;
	37540 : 1;
	37541 : 1;
	37542 : 1;
	37543 : 1;
	37544 : 1;
	37545 : 1;
	37546 : 1;
	37547 : 1;
	37548 : 1;
	37549 : 1;
	37550 : 1;
	37551 : 1;
	37552 : 1;
	37553 : 1;
	37554 : 1;
	37555 : 1;
	37556 : 1;
	37557 : 1;
	37558 : 1;
	37559 : 1;
	37560 : 1;
	37561 : 1;
	37562 : 1;
	37563 : 1;
	37564 : 1;
	37565 : 1;
	37566 : 1;
	37567 : 1;
	37568 : 1;
	37569 : 1;
	37570 : 1;
	37571 : 1;
	37572 : 1;
	37573 : 1;
	37574 : 1;
	37575 : 1;
	37576 : 1;
	37577 : 1;
	37578 : 1;
	37579 : 1;
	37580 : 1;
	37581 : 1;
	37582 : 1;
	37583 : 0;
	37584 : 1;
	37585 : 1;
	37586 : 1;
	37587 : 1;
	37588 : 1;
	37589 : 1;
	37590 : 1;
	37591 : 1;
	37592 : 1;
	37593 : 1;
	37594 : 1;
	37595 : 1;
	37596 : 1;
	37597 : 1;
	37598 : 1;
	37599 : 1;
	37600 : 1;
	37601 : 1;
	37602 : 1;
	37603 : 1;
	37604 : 1;
	37605 : 1;
	37606 : 1;
	37607 : 1;
	37608 : 1;
	37609 : 1;
	37610 : 1;
	37611 : 1;
	37612 : 1;
	37613 : 1;
	37614 : 1;
	37615 : 1;
	37616 : 1;
	37617 : 1;
	37618 : 1;
	37619 : 1;
	37620 : 1;
	37621 : 1;
	37622 : 1;
	37623 : 1;
	37624 : 1;
	37625 : 1;
	37626 : 1;
	37627 : 1;
	37628 : 1;
	37629 : 1;
	37630 : 1;
	37631 : 1;
	37632 : 1;
	37633 : 1;
	37634 : 1;
	37635 : 1;
	37636 : 1;
	37637 : 1;
	37638 : 1;
	37639 : 1;
	37640 : 1;
	37641 : 1;
	37642 : 1;
	37643 : 1;
	37644 : 1;
	37645 : 1;
	37646 : 1;
	37647 : 1;
	37648 : 1;
	37649 : 1;
	37650 : 0;
	37651 : 0;
	37652 : 0;
	37653 : 1;
	37654 : 1;
	37655 : 1;
	37656 : 1;
	37657 : 1;
	37658 : 1;
	37659 : 1;
	37660 : 1;
	37661 : 1;
	37662 : 0;
	37663 : 0;
	37664 : 1;
	37665 : 1;
	37666 : 1;
	37667 : 1;
	37668 : 1;
	37669 : 1;
	37670 : 1;
	37671 : 1;
	37672 : 1;
	37673 : 1;
	37674 : 1;
	37675 : 1;
	37676 : 1;
	37677 : 1;
	37678 : 1;
	37679 : 1;
	37680 : 1;
	37681 : 1;
	37682 : 1;
	37683 : 1;
	37684 : 1;
	37685 : 1;
	37686 : 1;
	37687 : 1;
	37688 : 1;
	37689 : 1;
	37690 : 1;
	37691 : 1;
	37692 : 1;
	37693 : 1;
	37694 : 1;
	37695 : 1;
	37696 : 1;
	37697 : 1;
	37698 : 1;
	37699 : 1;
	37700 : 1;
	37701 : 1;
	37702 : 1;
	37703 : 1;
	37704 : 1;
	37705 : 1;
	37706 : 1;
	37707 : 1;
	37708 : 1;
	37709 : 1;
	37710 : 1;
	37711 : 1;
	37712 : 1;
	37713 : 1;
	37714 : 1;
	37715 : 1;
	37716 : 1;
	37717 : 1;
	37718 : 1;
	37719 : 1;
	37720 : 1;
	37721 : 1;
	37722 : 1;
	37723 : 1;
	37724 : 1;
	37725 : 1;
	37726 : 1;
	37727 : 1;
	37728 : 1;
	37729 : 1;
	37730 : 1;
	37731 : 1;
	37732 : 1;
	37733 : 1;
	37734 : 1;
	37735 : 1;
	37736 : 1;
	37737 : 1;
	37738 : 1;
	37739 : 1;
	37740 : 1;
	37741 : 1;
	37742 : 1;
	37743 : 1;
	37744 : 1;
	37745 : 1;
	37746 : 1;
	37747 : 1;
	37748 : 1;
	37749 : 1;
	37750 : 1;
	37751 : 1;
	37752 : 1;
	37753 : 1;
	37754 : 1;
	37755 : 1;
	37756 : 1;
	37757 : 1;
	37758 : 1;
	37759 : 1;
	37760 : 1;
	37761 : 1;
	37762 : 1;
	37763 : 1;
	37764 : 1;
	37765 : 1;
	37766 : 1;
	37767 : 1;
	37768 : 1;
	37769 : 1;
	37770 : 1;
	37771 : 1;
	37772 : 1;
	37773 : 1;
	37774 : 1;
	37775 : 1;
	37776 : 1;
	37777 : 1;
	37778 : 1;
	37779 : 1;
	37780 : 1;
	37781 : 1;
	37782 : 1;
	37783 : 1;
	37784 : 1;
	37785 : 1;
	37786 : 1;
	37787 : 1;
	37788 : 1;
	37789 : 1;
	37790 : 1;
	37791 : 1;
	37792 : 1;
	37793 : 1;
	37794 : 1;
	37795 : 1;
	37796 : 1;
	37797 : 1;
	37798 : 1;
	37799 : 1;
	37800 : 1;
	37801 : 1;
	37802 : 1;
	37803 : 1;
	37804 : 1;
	37805 : 1;
	37806 : 1;
	37807 : 1;
	37808 : 1;
	37809 : 1;
	37810 : 1;
	37811 : 1;
	37812 : 1;
	37813 : 1;
	37814 : 1;
	37815 : 1;
	37816 : 1;
	37817 : 1;
	37818 : 1;
	37819 : 1;
	37820 : 1;
	37821 : 1;
	37822 : 1;
	37823 : 1;
	37824 : 1;
	37825 : 1;
	37826 : 1;
	37827 : 1;
	37828 : 1;
	37829 : 1;
	37830 : 1;
	37831 : 1;
	37832 : 1;
	37833 : 1;
	37834 : 1;
	37835 : 1;
	37836 : 1;
	37837 : 1;
	37838 : 1;
	37839 : 1;
	37840 : 1;
	37841 : 1;
	37842 : 1;
	37843 : 1;
	37844 : 1;
	37845 : 1;
	37846 : 1;
	37847 : 1;
	37848 : 1;
	37849 : 1;
	37850 : 1;
	37851 : 1;
	37852 : 1;
	37853 : 1;
	37854 : 1;
	37855 : 1;
	37856 : 1;
	37857 : 1;
	37858 : 1;
	37859 : 1;
	37860 : 1;
	37861 : 1;
	37862 : 1;
	37863 : 1;
	37864 : 1;
	37865 : 1;
	37866 : 1;
	37867 : 1;
	37868 : 1;
	37869 : 1;
	37870 : 1;
	37871 : 1;
	37872 : 1;
	37873 : 1;
	37874 : 1;
	37875 : 1;
	37876 : 1;
	37877 : 1;
	37878 : 1;
	37879 : 1;
	37880 : 1;
	37881 : 1;
	37882 : 1;
	37883 : 1;
	37884 : 1;
	37885 : 1;
	37886 : 1;
	37887 : 1;
	37888 : 1;
	37889 : 1;
	37890 : 1;
	37891 : 1;
	37892 : 1;
	37893 : 1;
	37894 : 1;
	37895 : 1;
	37896 : 1;
	37897 : 1;
	37898 : 1;
	37899 : 1;
	37900 : 1;
	37901 : 1;
	37902 : 1;
	37903 : 1;
	37904 : 1;
	37905 : 1;
	37906 : 1;
	37907 : 1;
	37908 : 1;
	37909 : 1;
	37910 : 1;
	37911 : 1;
	37912 : 1;
	37913 : 1;
	37914 : 1;
	37915 : 1;
	37916 : 1;
	37917 : 1;
	37918 : 1;
	37919 : 1;
	37920 : 1;
	37921 : 1;
	37922 : 1;
	37923 : 1;
	37924 : 1;
	37925 : 1;
	37926 : 1;
	37927 : 1;
	37928 : 1;
	37929 : 1;
	37930 : 1;
	37931 : 1;
	37932 : 1;
	37933 : 1;
	37934 : 1;
	37935 : 1;
	37936 : 1;
	37937 : 1;
	37938 : 1;
	37939 : 1;
	37940 : 1;
	37941 : 1;
	37942 : 1;
	37943 : 1;
	37944 : 1;
	37945 : 1;
	37946 : 1;
	37947 : 1;
	37948 : 1;
	37949 : 1;
	37950 : 1;
	37951 : 1;
	37952 : 1;
	37953 : 1;
	37954 : 1;
	37955 : 1;
	37956 : 1;
	37957 : 1;
	37958 : 1;
	37959 : 1;
	37960 : 1;
	37961 : 1;
	37962 : 1;
	37963 : 1;
	37964 : 1;
	37965 : 1;
	37966 : 1;
	37967 : 1;
	37968 : 1;
	37969 : 1;
	37970 : 1;
	37971 : 1;
	37972 : 1;
	37973 : 1;
	37974 : 1;
	37975 : 1;
	37976 : 1;
	37977 : 1;
	37978 : 1;
	37979 : 1;
	37980 : 1;
	37981 : 1;
	37982 : 1;
	37983 : 1;
	37984 : 1;
	37985 : 1;
	37986 : 1;
	37987 : 1;
	37988 : 1;
	37989 : 1;
	37990 : 1;
	37991 : 1;
	37992 : 1;
	37993 : 1;
	37994 : 1;
	37995 : 1;
	37996 : 1;
	37997 : 1;
	37998 : 1;
	37999 : 1;
	38000 : 1;
	38001 : 1;
	38002 : 1;
	38003 : 1;
	38004 : 1;
	38005 : 1;
	38006 : 1;
	38007 : 1;
	38008 : 1;
	38009 : 1;
	38010 : 1;
	38011 : 1;
	38012 : 1;
	38013 : 1;
	38014 : 1;
	38015 : 1;
	38016 : 1;
	38017 : 1;
	38018 : 1;
	38019 : 1;
	38020 : 1;
	38021 : 1;
	38022 : 1;
	38023 : 1;
	38024 : 1;
	38025 : 1;
	38026 : 1;
	38027 : 1;
	38028 : 1;
	38029 : 1;
	38030 : 1;
	38031 : 1;
	38032 : 1;
	38033 : 1;
	38034 : 1;
	38035 : 1;
	38036 : 1;
	38037 : 1;
	38038 : 1;
	38039 : 1;
	38040 : 1;
	38041 : 1;
	38042 : 1;
	38043 : 1;
	38044 : 1;
	38045 : 1;
	38046 : 1;
	38047 : 1;
	38048 : 1;
	38049 : 1;
	38050 : 1;
	38051 : 1;
	38052 : 1;
	38053 : 1;
	38054 : 1;
	38055 : 1;
	38056 : 1;
	38057 : 1;
	38058 : 1;
	38059 : 1;
	38060 : 1;
	38061 : 1;
	38062 : 1;
	38063 : 1;
	38064 : 1;
	38065 : 1;
	38066 : 1;
	38067 : 1;
	38068 : 1;
	38069 : 1;
	38070 : 1;
	38071 : 1;
	38072 : 1;
	38073 : 1;
	38074 : 1;
	38075 : 1;
	38076 : 1;
	38077 : 1;
	38078 : 1;
	38079 : 1;
	38080 : 1;
	38081 : 1;
	38082 : 1;
	38083 : 1;
	38084 : 1;
	38085 : 1;
	38086 : 1;
	38087 : 1;
	38088 : 1;
	38089 : 1;
	38090 : 1;
	38091 : 1;
	38092 : 1;
	38093 : 1;
	38094 : 1;
	38095 : 1;
	38096 : 1;
	38097 : 1;
	38098 : 1;
	38099 : 1;
	38100 : 1;
	38101 : 1;
	38102 : 1;
	38103 : 1;
	38104 : 1;
	38105 : 1;
	38106 : 1;
	38107 : 1;
	38108 : 1;
	38109 : 1;
	38110 : 1;
	38111 : 1;
	38112 : 1;
	38113 : 1;
	38114 : 1;
	38115 : 1;
	38116 : 1;
	38117 : 1;
	38118 : 1;
	38119 : 1;
	38120 : 1;
	38121 : 1;
	38122 : 1;
	38123 : 1;
	38124 : 1;
	38125 : 1;
	38126 : 1;
	38127 : 1;
	38128 : 1;
	38129 : 1;
	38130 : 1;
	38131 : 1;
	38132 : 1;
	38133 : 1;
	38134 : 1;
	38135 : 1;
	38136 : 1;
	38137 : 1;
	38138 : 1;
	38139 : 1;
	38140 : 1;
	38141 : 1;
	38142 : 1;
	38143 : 1;
	38144 : 1;
	38145 : 1;
	38146 : 1;
	38147 : 1;
	38148 : 1;
	38149 : 1;
	38150 : 1;
	38151 : 1;
	38152 : 1;
	38153 : 1;
	38154 : 1;
	38155 : 1;
	38156 : 1;
	38157 : 1;
	38158 : 1;
	38159 : 1;
	38160 : 1;
	38161 : 1;
	38162 : 1;
	38163 : 1;
	38164 : 1;
	38165 : 1;
	38166 : 1;
	38167 : 1;
	38168 : 1;
	38169 : 1;
	38170 : 1;
	38171 : 1;
	38172 : 1;
	38173 : 1;
	38174 : 1;
	38175 : 1;
	38176 : 1;
	38177 : 1;
	38178 : 1;
	38179 : 1;
	38180 : 1;
	38181 : 1;
	38182 : 1;
	38183 : 1;
	38184 : 1;
	38185 : 1;
	38186 : 1;
	38187 : 1;
	38188 : 1;
	38189 : 1;
	38190 : 1;
	38191 : 1;
	38192 : 1;
	38193 : 1;
	38194 : 1;
	38195 : 1;
	38196 : 1;
	38197 : 1;
	38198 : 1;
	38199 : 1;
	38200 : 1;
	38201 : 1;
	38202 : 1;
	38203 : 1;
	38204 : 1;
	38205 : 1;
	38206 : 1;
	38207 : 1;
	38208 : 1;
	38209 : 1;
	38210 : 1;
	38211 : 1;
	38212 : 1;
	38213 : 1;
	38214 : 1;
	38215 : 1;
	38216 : 1;
	38217 : 1;
	38218 : 1;
	38219 : 1;
	38220 : 1;
	38221 : 1;
	38222 : 1;
	38223 : 1;
	38224 : 1;
	38225 : 1;
	38226 : 1;
	38227 : 1;
	38228 : 1;
	38229 : 1;
	38230 : 1;
	38231 : 1;
	38232 : 1;
	38233 : 1;
	38234 : 1;
	38235 : 1;
	38236 : 1;
	38237 : 1;
	38238 : 1;
	38239 : 1;
	38240 : 1;
	38241 : 1;
	38242 : 1;
	38243 : 1;
	38244 : 1;
	38245 : 1;
	38246 : 1;
	38247 : 1;
	38248 : 1;
	38249 : 1;
	38250 : 1;
	38251 : 1;
	38252 : 1;
	38253 : 1;
	38254 : 1;
	38255 : 1;
	38256 : 1;
	38257 : 1;
	38258 : 1;
	38259 : 1;
	38260 : 1;
	38261 : 1;
	38262 : 1;
	38263 : 1;
	38264 : 1;
	38265 : 1;
	38266 : 1;
	38267 : 1;
	38268 : 1;
	38269 : 1;
	38270 : 1;
	38271 : 1;
	38272 : 1;
	38273 : 1;
	38274 : 1;
	38275 : 1;
	38276 : 1;
	38277 : 1;
	38278 : 1;
	38279 : 1;
	38280 : 1;
	38281 : 1;
	38282 : 1;
	38283 : 1;
	38284 : 1;
	38285 : 1;
	38286 : 1;
	38287 : 1;
	38288 : 1;
	38289 : 1;
	38290 : 1;
	38291 : 1;
	38292 : 1;
	38293 : 1;
	38294 : 1;
	38295 : 1;
	38296 : 1;
	38297 : 1;
	38298 : 1;
	38299 : 1;
	38300 : 1;
	38301 : 1;
	38302 : 1;
	38303 : 1;
	38304 : 1;
	38305 : 1;
	38306 : 1;
	38307 : 1;
	38308 : 1;
	38309 : 1;
	38310 : 1;
	38311 : 1;
	38312 : 1;
	38313 : 1;
	38314 : 1;
	38315 : 1;
	38316 : 1;
	38317 : 1;
	38318 : 1;
	38319 : 1;
	38320 : 1;
	38321 : 1;
	38322 : 1;
	38323 : 1;
	38324 : 1;
	38325 : 1;
	38326 : 1;
	38327 : 1;
	38328 : 1;
	38329 : 1;
	38330 : 1;
	38331 : 1;
	38332 : 1;
	38333 : 1;
	38334 : 1;
	38335 : 1;
	38336 : 1;
	38337 : 1;
	38338 : 1;
	38339 : 1;
	38340 : 1;
	38341 : 1;
	38342 : 1;
	38343 : 1;
	38344 : 1;
	38345 : 1;
	38346 : 1;
	38347 : 1;
	38348 : 1;
	38349 : 1;
	38350 : 1;
	38351 : 1;
	38352 : 1;
	38353 : 1;
	38354 : 1;
	38355 : 1;
	38356 : 1;
	38357 : 1;
	38358 : 1;
	38359 : 1;
	38360 : 1;
	38361 : 1;
	38362 : 1;
	38363 : 1;
	38364 : 1;
	38365 : 1;
	38366 : 1;
	38367 : 1;
	38368 : 1;
	38369 : 1;
	38370 : 1;
	38371 : 1;
	38372 : 1;
	38373 : 1;
	38374 : 1;
	38375 : 1;
	38376 : 1;
	38377 : 1;
	38378 : 1;
	38379 : 1;
	38380 : 1;
	38381 : 1;
	38382 : 1;
	38383 : 1;
	38384 : 1;
	38385 : 1;
	38386 : 1;
	38387 : 1;
	38388 : 1;
	38389 : 1;
	38390 : 1;
	38391 : 1;
	38392 : 1;
	38393 : 1;
	38394 : 1;
	38395 : 1;
	38396 : 1;
	38397 : 1;
	38398 : 1;
	38399 : 1;
    default : 1'b0;
endcase
end


endmodule