module control (input logic Clk, Run, Reset_Load_Clear
                output logic Clr_Ld, Shift, Add, Sub ) 

endmodule