module sext() //dk if we need to use
    #(parameter width = 8)
    (input logic [width])

endmodule